��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���麍�Ks�%$����+d7��/��������ߔ,���<�E�]��&��z>��>�X�����A�
&CʁRR���o>���q+�AR��k�b� B�����C(D�x)�d�!gN&{����+&f���^��T�JЬJ	yh�ldڪ��:RV۽�أv��椏����7�5G��Ξ@��/6����=;+�Cgt�ܫ����ߥo��yqa�ĝ!�G�F#{5� �E؃��\il����A�E�sƸ��]��i��Y���i���	��'i�6�9U�x� ��n���}FA3�[�����Pٵ&�����''�qe�-�?
�%w$�W��[��m�w�xH�O�I�	�@����[oVʭM�A��t��B�gx�K���8C��G#h�̾cZ���8���L1�}�L�RZ��L/��W�p���;lB��*�Y��4�%]�Y�:�b�\Yv_f��!P�{
2G�-�Pi���xhB�ё�&���7`��G%����U�^�9���t�M� ���X3���#���u�鉾μr|Wh��h��Kɟ������cG:��9J>:���ϔ"��nE��2�����>pS4s��	�(G4{(S�L�:U�.@�|R0�L8������j��IB�"���N������ys��ė/,ҊN	q�v�Z��\R�w�0xtʎ5x5�������v�7\M�k���%n;c-<�<;�`.���B1�7���[�D�\�A��fIj�)����懋�f�7`_�%�E�i�j��yF���^�s�[wg`}vёp�M�=&d.�ȩ$7l	�$����>&R=�M� N=;5k�B���t��7�@>j�c�� �����<�T�3���:����� ��	'
o 	�����v�E0=�(=S� �:$su��
�T��퐣�nXq�u0�pG%�κ6�t$k�%�,�er���p�����w��6���@����jV8U����3~ݦ�G�nM��D������g���擉}�0��j�j�������{2�p�L�i�׿�N��Զ+�H����C1A�*�j�P?��섇�"n��DVJ���9Յ`�Ľy�����.#[׋�2:^+{`�p�v�2�T��=Pi��H�<d�ȿ˖����}LL4�z��n�S2�>o�7����HK�/v'�]�HG�h+s	L�&�!&�B�C7qux����|M�e��q!|�v�M���5W��]��%=�ӥם��㭼�V�ֻ�����L\��,������,�a ��� ���)����k@��nד���|P ÿ���7kh�,.]
�/���n�2y�r��S�y����`E3Ct�ڤ�������&�[�*}���\ �4K6���)��~A�����|��H-x�F��*�V͙��E�x���Z�y�=�
�'�+���@{����f����EV���Θ8M�@*�R��4�d*:����+�~��z)s�c������~ i0�8b���[�f��{a R�2�M1��y�.Xq�A ���f!�x����}�}��n������Yf¼S����Ht�Ozŀ�p*��4����CD�`�+�l�9I�k_�̖u���P��X��K�q�EŨ�,J�����Bk�m�@̶t��IC�v؝��j���wH������&g�AQ��UHy�~�]�## G;U����Q���d���;(�f�~�����Ŵ3�5<�S\f�K
	Xaܶڰ���I��1L6�}�2@�����g-.��oV�0T6x$��u�����p����$�i���%c�uX��ُ6���������<��m�{�)��]�Ɛ���j}")�6x4E쿽�j�D�-�\�M1��r,�mT��Mq���D�i�n�3,IOf��pt�i��!RY92r��B�M�BV�hY@�����,�+��G�.Y�]}���G�	/��9���0�&�Q��H�E���U�ʺ*0������_�}V��]���P|�0�YLj��ci�"��3�w�
�$`�;������ ��U�z���ͱTo�\�o���M֫��DGf�q�}r�M�˔/��v,�y�`gt�y�iR��֢���G����J�f�#����Ls�n��g�(l�"�+��� zA���V�+d��O��	�H���!;]��[Z��J�7c���1����n2]��v�>1e�����r��iI_3�`a��� �@��u�����W����?pn�M�,S�#-U.���������'B��^P\\&����^�!'>3��H�,�HPƙ�+�tE	S�"{�+l+Q���`��4�dҿʛ�S�|� %�^C�7�x���`�;n#�u��W�p���Cd�QPF�5ܚ8=��V�����iN?}��m ���l��\���*�1���B^8�3���߉�h�P�S�����5��e�g�� ��<��H��\�x��y&�զ��e1��6�%�B�xL��U`�d��^��oړ�d N��\,B���V=��|kO�g"��0 i����0o�~ˑTG��@�(�����_����DG�eR%���^�uEn���BN��������<t����n�jEmgng��������;��p�5�(�e�T_�dƥ���!��}�5]�v%���??VL�cw�w���-#��'�>�]*�i�	�-�̪crN���׋�928�RRf�8���ks�uR���螰o����oﲚ��J�G������^��K�t����蚼��nWi�Q��.�#\�1����E$��JQ:\�f����cӬ����@n���i������ƶA�@�*7v�|�E^>�w�Z��r�tbF���z���n��J���8ܝ`\r5��Y��ą/��v`8��9�,AԬ��zZ�?O���oU���E����(�^��I~U�69캥�6��EM�9U+>*��)�I �h��,���q�Z!��Ͳ?����W��/@��
���4Ig�¨�p~t�v��W���1�n�
��& =��Če�۬+���*��}����"���n-p���ӠJ�O�Lo�ҝ��������P,�(E��������M�a�X�$��!���<&�����u�z9N����PKO�����3��h�窻l���Ƽ깁�S�Z08�q�;8LRy�F�^�m���/\;�����9χ^��)<v+(?��4������Kr�Lȸl:v%@X6P%c(�]9�V)`s;BOؽ:�,<�=E��%7�{��������K�vFYk�A��$��H�I}�Y�6>D9�Хn}�����a2KK�%�=UC۝����UV{,M��'������gꉻ��*�Z�5��ԥ����� �`7?��S�M�ܢw���{���26,�@I03�*h����ȇm�����ax�r�Y��C�X䭑'(pa�H��݆9݋�,[�,~%����@؝������(�o��!��X��d�G�=÷�\��S�ꝲ����}��{��B��N}IG��ށ��}��
�,�u���|���E�C����K��mM�ȇ9�^�HG��;��YKm���l�g��͒�L~��+^�N2�u�*�|�o�0��. ���V����:Z&�dcs�N��o�ݾ�|�D���\�d��]ΪS7t����)�ߕ���}�k#�:��
��(�R�}`^�����q/(��0hѳ�H�m��
@!�9l�?\�=�.��%��I�aw�����2&@��g,�~ܸ�?YQ�,�>H�ϣy���@�et�����b�M�i�����͹�w�⚄�ND�!+R	e����O�w��r������`����fL�F���w��w��/b˂U3ކ�=����r�BK`��w�bJL��#��q��񒴂����$Gps��yp��Go���,�@
H�����[k�z�j ��e�s����\%�"N9ws�<���ٓ
�l�կF��
Kh������j��X��G�W0�ZA��5)��P
7�T�Z��:��p<	�J��yњlj��b1�9s�[�I��*\���LxR�ј�Ʃ�WSy׊��o�6�+��份�U� %���|�{�Q{W�.��Q7���#rO���]��9�q�樲Ը΢��뫧.���.�=r��̓��@�ű�־������\�ibpר�7�W�P��%TDCّv���l[���q׼I$U�tK׮�ߩ�%��4B��^ �?%�ƅ
]�%�f<�(�|�H��`���!*݋�栳
�r���|�P2,W.�z���K~��%�h9�\�=8*��xQ],>(�b٭��l�
�`�6�(D4(`
׳�U����o<h�,���Ͳy�/$�T�Ѫ]���s��&���52R�[�A���J����3Hf{n�?:s�х���������2�5�>ɞ���j*t�̷Ra!5l�*�-p�Ӹ =Z��VV�p4��A�7��0����P2/
��/j���������mܝ.{�:&�� ��3�3��O
GVU,�rn� �Y�P���(q��b�)q%O�0�do���;�_?�r4�Х �y��M�%A}���ۈT��mi��e��*F�5��π�>���SL��K3���5�l��J�L�����E3W�˗�>��;dX�<��*�v;����k8ī�`�DN���N��l�������I�V#?����bM�5U���$�(���x	�]�;D�x�Df|Bg� >_Q�a'Ͽ�h��<�	L�����ՃL�u� h�br��O�ķ%� ~8�u/E�S9�պΩ+]�y��+��ӵ����&)@��W���2�"��V���-���Q���u�Ą�����u�Ɯ���v��tW�8+W�!"�p��p��~.���9�}����ѫB���m��W^MX����x��q�9ݱ���?ZG;� ��aUy���R�eD3���a��s0�6Z��k�i�,����"֤� ֘�1?�g�)���|��jW@5ߟ�Җzٸ�ӿ��)E&s��0W���p�~�'�/ʯǚ���սΗZD�
'Xy�u��1��N��Bg&�7m��dp+E���@�A �5B�a�b���N���t�	8ԫ�n�>��DI��!y�	�<�Q)�%�;��H���t�F1��d@��F���>���ѯ��%�neY�����HBG���N����b�A8J�T�`j���n�4X��������M�pV�.��]�<���=Bw$��k�O�������yIH�eUE�j�i�luR!B�Х�����eZ�I�;S:6c-��/��lBL�X)L�j�$�(Aψ�&
)�_���D;�i��v�oH�T��l֚��#��-���*>�Bh�1�����b�-!\p����hW.D��Y���wu"a�-؊�Ҳn2gA���&!/;�\�	�|TW��q�X�t��Z�P��(y���$É�;_0�bjƺ�*�ɓ�aG��M���Pٹ5�o�iDvx���1���5j���?�.ﰈ�����'�O2�d�?�uQj� %�i��9C�J{�UR
ӣ	'����G�VC�m�q{x+-�X~s����}�bPK���E���T�ࡖ�>ojgX����"\2o�nb��%@?>g�|����<���\c!��ʐ�;䲁b��k�X�fh��C��j3n�dTxFR�B�mr��?ix�D*���c��"�^���Y	�x�wf~s-�Ra�&��c��#r�iK[���j������!{rkt��b6zB�����2jt��9Q�[��;���?�T;եMYx�8���1�A����Ǡ�$�;�Qh������n��A�t6	6��z�i�ˊ�")iI�*nT�28,��);�4M����*��p�hޤ�آ�M����+��X��X����D��˨+�_��+�N_e�����ԾI��4�.�z�|��7�v,�e�?�X���J�w/�`�Q��v��6KW�H��=[RCZ��d�M"BY�G����!Z�Kv	1��8y�0��+'���^eH�NZ��/����/y�V�O���>���	��&9u���\��J������xYC�: N�T��"��2����AF2ro�N�F/������洽Ͻ�Ŏ�⢃�m��5��W�� ��x�q�8D��Ģȣ��l�h:]�bw��	����T=c��K^�x�Ɵ�x:��j�^uG���N��n�xF
ս�z�h]b�$��p)�x
Z�aŬ�:��0r�*.����L�f9:c���Dpi��_�G /��Z�4���[+���-�Y�����=����9b�+��W���@g:��֮����w1s3M'�I��VhD�lGe�qOH�g��.�v�O9��bj��a�T�sEU#���\�i�˝W���/�Ý�+n���0�V����.�]��(�&{"�l*���Z۲��??(�wDCj5�l)w�N������[jл�5�NS}��ȅ7�E�`J�4��� �"���|Y��/�^��������)n���vy���ʶ8kܝ�])��x��{mth7��&���4%��5M���C��z޲��Bv��7�+ɤ�>�B��8����'H��E}���mz�p��~^LB�m��NH.`oMw����Yo~�zK��tdӟ�Ew��7���o�7?U�٥0�I����.���ݘ�$�v��z����J��e-����Ð�qR��ɗ�%�B�o�RY�,�u�$��h�\I2f��z��Aܯt˕ ���$M@T�?6u�z?�G��t�.�c������}+b����a��<�%����Il�3#cs>T��ʚ��M
�`���7��*�w�A�O�=�h4���O�J;~Ο$�ĤN�����U�=��k�X�q�I@9 �a�&ث�S�T���ʛU�k��έ�t� 
�s�a_�
��Zy��{&�j����}��jS����"��v�CW�{ḍ�"�����H��3�8/���1���*���,���$ɪϽ���Y�#�L��K	��f纽7�i���P�ǂ��t����:��G�o�+Q(˸���y^4�m���IYp�����O*���F��M��S��jz*ml��ȒEz�i����{�^�$ۆaS*[.Q�)�ḁi�v�W�rτ+����)�!�W+��k�� ��f�[v�zb�0�2B���p'T?�q����.�\D��Q�Eχ�Y��G-��ƨ�~ub��D�÷*|X���~Uo�HI�"��gh5}!NY�d��o���5��q���/�Y-�".^9�u?5e��\�J:�(��%�iˢU���,Z��eZ�h���*7@�F�6��3�q���=G�*V �߀ȕ�����z'!���6�Ƒ��ͫ��cB�>.��]��o����YIs��|L�.��B���m�,�DP��������*oi�5���]���~���
}$���$u��T�p��Cw��[��@�k��課��q���+΅QV��U�H��I�Ul<��W��"�%io_��f����AjS�Sp�b�5;��b��0MQ�p���٦z6k�L�#=qi�^���1Mw޻�D��:ͣ�tmrR��Հ�'�͔C��	%��l�.�O�,#8g���ך�v���+��w�U'kʖ@�������GX��x^4?���^��T�V���_�GV�Qc�ء�=��nn���k�( �c�yiNQ�����pl��eGz��l�Ԃ���?:���-D��eu2��:P�(y4��Eη��¾4�����~�&V\Gܰ�|�+��	09y��lr�ã�+��;�:f�jܭ�:K>!=@���;�>�{����ِL~R��d����ʂ9�Z>f�!�^g����^WF��^�-��bhR��8ZC"�a~�Z?X"�h����.�a/6K�߽�P�k������:k0�0�5O���XQ+�w̡k�'�H)�e�Rě��b�~�pq�f��,��&��(<x�>"�HXت����Y�E��� _f�u%�bTv�W/��Iq�Ŏ)b����N��
o&���?!W�y̳���� �O��ܑL���i��F2bN�[�����-��.%�)Ƞϫm�#ϟ�_��@1�������$���ڳ~��;0�����ۮ��=�*`��#Q��?��f�c�؍q�e<�?A����J����}� ̪
�;�Fn�|I�4'�L-yF[E�,�H:z2���������xp�q�|Bt뚿��.��b���d�eWb��O��1��(�e���tK����lHa��Ӈp��d��jq�!�3�4�H�k6~�~9�%�|��k�]{�?�m�ڍ��^W�l�gԶDEU���o��[ڽ�x����P�n���{h8�:s[w�d{���:�,���g,�P䜄��5�{�Ka����t�s� � 
9�>������@ģ)��`��绞[����d��LvH�h�+����v7�H����B��A������]���5AрL�Q�1�t+���=��;2U�5w!�f�?�/�h=B�.�;��˸$x���kh�xnG�jMe�CTQU�V"�x��ж<��hP�d�/'9�q���?7С���PI�-ʴ<~�rz�I���pPs�i	t��>`���xVT�x݃�Ft�NA��ܠo���P3�hix,BŞ��lhֽ��r�h�G�T-Vpc�с��=�
�E� 6Z�u��x	47,A�.\�-`¦x���/^XR��4�ߺ�=�>ɹT�{�²��|���� �8�:����W"�]�t>A��8!����ʔ�WH�"Nu��d��l��A���>�[���,g���0����6cٛaI�}֧Jז=y��F]��o�rq�%J�^F1=�8
Na6������ ̯��^���%�Mז"�Xm�A��._�ů4��6�!wY�oD���ꊋ�m�(M�3�3ϱ S>�T���V���S��R/s_"K"��������vG�k`>僀�<���������ikl������#�9��ȝ8͵~w� �|e����8�d�.�-�q_U��g���V��rS�O�V|V  X�A���4()Ĕ�`�ף6-}�,�S�UG��ĶB�نn��P��>EK�t�w4�"�[�Y����S�?eB�+"���gܥ!	��R���3~1R��{Ps٢;9{سSٰ�7tzF'�ܶ��Iŀ�5�w!�E�|�9��$S��	�z?ͱšz�|V��ᝎ�<B){�!�?�O�G� �`-�<���z	��lF���o�LG��Vqiq�����Q����5j�M��Π>���?�HGXe�||��5͇߂�7���lE,}��� �Y8�g�ʤn�+����3�����{0B©�YɊ˶�����b�a݆
��#��H-M��i��e��� �@I����2��]���xoD���׽S鳬LB�+��TNnQ�����?	ѽ��R<1�Ez�p�щ�7�������k��k+1F��mw�:�a�Il�3�B�W��`̢���y�T�E�.|��O�j˞��ޢ�"�K��?1u�����&z{\u=�w�s�!���Y�&��sV�٤7 ꡕ��ӟ�MS|���\�ҝ��씇�����>"�TOf�?_R��Ac�0�
�ox��?11f�R2�E"-�3N��y.X�@�����Օ��}���+�3vZ���筣rG����әA��Ҟ�O�ھ��4��)�*N٘�>Ңz�iG��O��u)����AF�\�Η�-��(Lƛ�ts,,�?��W
\���I������q�6Ԓn;F�ƞB%�����bn�p�W��H�w�s�A�;�R�n7N]Jɛ[c�?.�o�w&6~L�:���`�E�zq�r����O�l�S�ݝ�'��<B�f\9ga:�a!�'�5�_�GȬ:�}����O�>���o�����A���|=��ym�4���h�AG2z�O/��&�O7��_n\��AN/|�22e}�&щz�'Ҳ�k���`8����d�x6��q`le��3���췶|[�79����
�Q�J��N�[)�g�_$6=n��rl������Uً�6*{	��v�Q�:�N�!3O�E��OK��J�U�;����u�]l���zQX�iv�c�h�,�ut���"F[�.!@v����A���^V ���<|��:v�7�_4X �%C���l���)m�����ժ��u�c���������?��Ҥx�-�]��J��KL,�$��O�z�x��E]��C�/)|��j�Uhj��r��%S�k�t����c��q0�w��A1[��X:�ѫ�
g{#�2�J�\^���>�Z�<�#\����h��Ώ�r�M}$j��:n��}?�l��͇��r��s�\�(�F%�7y{���?�Q�ϣɑ[��M�oK܃CBj��k�5�!9[�����x�Q�e����V"�BeiÏ����v�dhC�.�jN��oЊ8�+s��^��%�HH�{	RW����0�c�L��(�c�α%��o@�R�U�K�2� T�h��\;q���X$.�G	?����a��-��1ȟA]L�c��>��b��k�f�/��)D���	ܵ7gT�0�
�*:����R�pU�S�1�0ӵ��3܇\�����W+�gp?�z�GZ�]ڟW�Ǒ/#`Cq���Dm2]�q�Ѕ,����o�Y! $JrO*�,B@KLl=U�	3�8��
�c�8bw��i6�Y������=��a��^��qB���[�o:��u�<�@Jդ�1krnt�LO�p��:u�3���Boc��+�$���$�/
n@�����QT9gW巒�Ǔ=k�s�T&A�U��g�=7�V�2��()1�`VРbR�k�����=�U��y�.����أ>3���c3� �T�n�gQP�[��-qYf�D�|�'���5��𜠴GE�wk�]>�C�v>���.�j�� ����A��*%*��㭟=�����S��-"Eế�!��# _	DUtv�<mTn�l�Z�U,�]o�/�
���Fz�c�I�!�*�EI�R[�{Q�� '@D�O� �d���d�u;�̇)YK��=�s�P#NXH6�SL�9P�]r����FdQ�0O}�r���<L*������ʓ�S�*� ��/��F���j���j���$H�MJ� *�~�e���c�$�ņd�E�ҎT�O��pz�"uO|�)z�����m_��G�����M~�r�`)�i�$�̓�Z	ӆ0�е�����L�U��#��Y3�y��_��HZj��J%8�3!I��k��3�fX�_�0ʹ$��c�%���V�_���`?��+32�X��r`��|x"�:=�_Տ#��l�bnս�w0���	�q��^�4��{}6�}���.����5^�	�Qj�v{YFAym;"h@�J�^�i�pF��a�W�`���:czB^e����1�CdK#�I��L���g���H�f��˹fwx��.��Lyɧ��gg����سY�a��k���m��~�Q�ć�p��W�=%zԟ��
���3�Tn]QYڢ_&�;���V�?�(�۾�D
U���;*w\�/���7QoU����H�g�� �zS����+��p�z��/�6 ��L���*�l�]$f�"~yPB������c�Y'�o�5�۵��
۪��c5�S���P�sU�_,��E�6����_>ѾM�[b��@n����P6�!��Z_�$,m��U��S����V��!c��$T��g�ZE��1��2)�'t��6�0�N�o��։ɓ��%o����b�?�`��|�(ֆ�B	���OZ'�)������A�MGK��rj&�3�G���W��-�C�YMQ��3�G
Wq"���Mc�qڝ�H,'�XWrf���*���d�h�x� � ����檇�����kw�6 ���A6x�vV���1�󃚰@�S#�e�t}>�Qr������Ai.��b-`��J��K� ��-�ҫ�o��7�ނ��n�jP�,F�h�����`�O�	��"��������)�S���0�A6�A�m���Iu5�ǥXjpn��5�>��R����\vS��^m7�I��ߒX���ϐl=UW>X���C�H��?�'$7����W����)��׍gu �Qٟ��H3�UJ���-y_6Z�0��V�g�^�K�n�\�0�� ��;��OЍMZCV�]6�]��$j����ʣ��+�"�u��[u�{��~��t��&���"���DM��6���bH�][���mS�q4''X~?��6x��?�Y;yڴs�)�����*(�*.��'"�#6�jsO{��r�D�:L׫pl�-�tl *rL����A�`㗢$Ń�VCG�t����~�3|�����S_"g�A78?0����˱)9?���Kl���5�L��:�Ap�(�d! �L
�a�M`x�5�2�<���n�6�G�H���[p�̄	7aVyv���.��t1�P��n�f>S�2��s��Z&F&� �;�IA��CҞ���䂛�ӭ�_�]+���r*{� �'���:�s5R$@Ԋ*�����k��L:�N�P�f�� �|��_�& ����';����C��Y/�C}��}'e��:���s�ྩ�޾��Z�4�9+AL��󑬸�L�ob����,v/[�I��*��BPE�y���=��#s���"$�½#��%��a�G�oKȨ��|ܴ�@��l�fF��^����,^����q���}��֛%| ���V�o<�yL�8�7�&)F�o-��Y�+���g��{�l]���J8�Bw���!���S�û��9�0�r�^�
Xs
��ϙ�����l�W�6�z.ǆ��h㩮X�$�_��`x�n$(.7!�:�^�A�3L����I�4��^ad��>�(�A�c�)=ռ�q�C�;<�'�������ӟn>Tҙm�>�x`���X&h*�/S�?Խn
{{esa�w�W���d�0�0yҷ}���8�3�f�d߄�c�,� ��p��uB �U������B�o�L�Z��9��P���(E��+�O�b�{��F0���y)�K���0`�n`���cHB��3�v��E�����~���zJur�cU�0wv���he�+=�4���ɩC���W>=��;.\g�ť�AD����		��wf_x�p1�(Ā!���e�q1	�U�,����`��_[m���	R.�~_�[9��O��F|�1�#"C�c�Z�[� �����B]u�3�[�q��|*�w�;s~x�p���^"CX /L�T�p�9�U:%K�b]6p�!t�{^��W�B�+Ԙ��'@��C�	*w.�*�%�z�{�0cQ;1ly���{��#Y5�L�/�-��������z�S�0�2�H�%րذb�"���7�zeE�����e�-�M���nF��m�~ݓd�쭭�9���� �TTgԜh���P�-N�zOqv�&�B����$�Ő�c�n�22Nݷ�=�<:�M�^�t�>�c�ȧ4�*�;�m�r��imu�+��
HL�}Hwՙ���g��j羳����~�֯ ��Ά������4zg�@ƪj�L�0�rW�y$k7I��MƼOԲ�ñ�h^�d$`�\�l��y�Vuz ��T==��V޲����ݿ[L�XH����+<���ݨ���uﰯ��7�}b������竴e�+����, ��z�HN{��#l��͌���#v�:Q�`bГ��.�����:���1��7AoχF;d��Z[����skVl�p�p��+�Ox����i��n�V�!t>�g����널O
�C�jW�B_�=r:�l��_��eI�p��~�[Q?K6�j<}a��]
/ũ=9L2>`�)K)W��Vn�� 	�`K�Y;������Z��Q6�:z_1��B�~�~3Z"�/5d��;b��\Naʵ�׵J�I�YQ��}z���b�6��o�X\�S�Cp���u�ʵ�S��gS�GZzvх���w��<����r�$��+E��& ~���
�<45�����e��a�i�,�v���/D�-��f���l&0rf�xw�E�f�ˏx�O��;J�(�?6d�r����/���i�����b���|��`?T���S �T^���D�pxiY�Y�""�6��T}:��Zf3`$i-�'4�+jKY/~0~H	���gIʂ�u)\�X �O�-'��I�5B�;J0`��[�q<%�v�+���d�32��@IS
���ekz�&�O��Г0�[�%�;)�E�	0꒿�\�\��"y2�	�Z!/Zq%��9� ���|m�00�Z�ä�m����ͅ���<?`����u�:��=&q6	�>��6��{G�Gc����T��}�v���,���EMj�)��Bu����ڭ� ;�����~x4t�_Uq^�����N3�yc�jf��@D��3�x�:�d�'�
c�%����e�K}|O�\�t�~�	j���.�ݬ�\�����0[��ܟd4n�W��w�[<��}��+�I j�����3���X��ɘ�ӳ(�/P�Y��T��΄q�e����0�ɫ�2p9&�߼�g�SQ0��-:��o�U.ߗ)?��썜0��;yԨ
��F��*���b��7X�������j���<�%��EK۫@�EE	��>�T��U_��J�X4�y��A��K]S�s	���)��I�8��������\D�p2���3�0��c����p�m��AG�z�$�Պv�:���vkv���m�-ڋ��1��n�B{b���@^՜v��>}Ŀ8���x�;X��v8��v�X���mo���ah���9�S3fM�EZ�N`�0-n���#��ċݺ���z���b
����#$����|±Q~��1�(�r�J0͟���`�[�F�0�s}��t��n6+ƴ
r�[��^�0@$�[��W�ӑ�@6�_�~M��3�꾣�1�w[k�ӵd+1�K��&���YM;��N���nޗf�+���ޯY5��tPMa�m&�#�w Q+.E;d���Pg��<��|0פ+�F�:���b;��=�{��Av������@X�R%t�~�%]��?cU���ʭZ�hjGg���r�u���*��3֝�����/	jP*�"�KV��� C��R�|�e,BnLoH��Cu����W���*󙆥o��:^�X�p��A�ks�}{%P�G����@/����1z=N���u|z{'��,b�m�x�8����ou�C��I��[�I��]Ee�2\r�u}@6��q
�.b���#���,痠C`T�'��s�'�!e"���� $���"���)����IR-�Dھ1�>m�H-���'�0�m7]�1�LطxJ�T1C��NC�/�WҪlEX���Z�i��͖�t����L���V��n׼�D�a���^G(4r�[��7!�l��9��"CQ�d0Q�N<'�鲈jj��_�s����p6�����,�<�L�j�
55#���'?N:5����������&�{��B;�>�
!��o��<���_�"�y�B+D�Ux�x��X��xR{�	�OD��7�SJ%UF�+�o�2u��vqE}ػ��pɦ<B�u�G6�|��kH&Q;�?���%�9K67������6�F\'y�Z��g$oe�� t�WՅ���(���@W��"��
x��`uQd���Νüy�����p����Z�"�wQ�g�yw�$�Q�ZR�L�pT�K����M֦q�[I���@Bo��B�0�F���Q߯�����/;V:�������4��o�ER��]�an���D�ŪOԽ�.�1��C�f,u+�]��p�/��"��q�?Q�s����݇�������β��˸ֿj?��(��O�>K��x��5¾�C]�eH��n�(;��xp�b�ų����踃��*gɣj
����n�"=�KQir�J&�P�^}��D�S��牼�m������K���G���2�Cr'J|Cf�I���aԖ2�47"6��EG8��:��{Ҟ�OH���f @?��H��7F$d�w�	o���m?�H0���5>jVR���;��^e�*H\Rq�"xhgCgb����-��fQ���rA�n�q=�I@�����8Z���|�/PW�P%�l����w�7�Qp��#��UI��)b���u�aB%U��+��$[H���6�����vb��uk6�ɴlr�+?�[0Um�an����qԩM����_��VeD�b=�ދ޿�)�����2qK���΄t^;��(dfu�8���{�qe׼�����$f~:�9�4�k)םX�5�$&$�ö���y�Ȥ&8`�L����^#�����t�v���/�Y��[����*�^�4�����?$��U;�jl���!A�?܏���c-�PM� �9G��M`�ּTe{���.�١Q��`O�>֏�s���=�\!�]D�Z:�H�G��@o��s��ƌ��u����x�}Ƚ�֌W�/G�U�'�L���RW2	u�h���|Ϥ�d�|YԚ�AdtC�b��٘��e��&��/z�
L��$k,����h3�襱���
��8�,	:]-���]�S�z����o,;/�ň,sr�f��N+C��w'���_�33{�Li�����
�6�%~�2 �͆�/e[��;G�a�t �}|(�.�3�Z'�4�m�]�Wd�t��-�MY��b��p�K�6��v�z�=TW�x��Vw���/�6�!OI�-e�j3�������˛`��K��U�Ç�%��ځ��Х(_-}�v�c��LJ;�1��Ru�x�RL�����I���x���K��Ij�s(֧Ik�gy�4~3h0f��E���%|,���W�NC��� {�y_��+1^@*!%/���a�1�s^�d�S���W�IY�J�|#G�IO��Ĥ�-Ra-11Eӊ��7wp�G܋�����X�g�Hxr��Bd�l� Cc��CЦi����Pq7��^��@��3��������UzYc^��e$h.�}s�ɑ~�-u�p&i+�![�\o�H7��x�3f�B�8ߨ�p���t�[��S��#>�c/{K�?<�pU����K`�vb�ƿo�&\)���عs�n��<��Q���N^���;�d���-e���P�sw԰ 黶23���<�ϴ����q!:��� � J�M�\p+.��l�^֠���q�iBG~$&��4q0|�I6V�ʍ����o���ؤ�th�m��Ҍ�����@��'m�5�q�_�8%�S#;2�dV��w��*�,6GZsa�ȁx�}/��~�o<�M�#Fd1����2�`��0��8�1�5R���͜y����>���x�&v�?^?E��~�(	?�.�M�ڡ�gHTB����ԣ&�ỊvBg58Z rQj�]�������n����BM�DYC���y>����8�+�4k�K����lߦ[;�/���c��� �O�Z?�t��^��c�Xri���%��!�}bB��'~LI|x�hP��@��?
��D �?�F��5I|N� K�WcLy%Zy��2�QOK�R����fh3n0��tqX�^l1*ɺ��I�$�?c6f�"�1����mA&�ߜ�Eh��{f�I.\�p�A�c[W��1ti��E֗5�z�J�X1~��pO��|֙qW\2���)��C��E����N;����É�I�uF�^��$JUP�6��P�B���|?�3�1s K���(k^���{/���&�2��������S@�.�T��"�s�FF�p���m�'q��F^9��^?i��_�C���KTS7�$
"YU�ښGY�0��ܷ���X���J��Ȁ��k����o��eK��t�G� ��]m�a�#���|.�I�{l۲���;�&Vfjr���*H1�����&&0Ded�]pB�51�#��f�$�ݧ�1���P�e9�*�򈍣2Tj��F�A��FP[�6Cdtc�z ���oLU�k�������_�$��P��b��rRW�!�R�@ez�t�5�=a��&WI>s
�̏1t�,	��C!~X����	������/ѱKuF�*g}��^\a�^L���WM����y����>YE��44���N�*�Ů���}��lo7؞I�딼s"6	n�ʛ:3�/��
ט^�H��+gAy�5� {��43L��3�S��j���_U��m�Pk��~��������I��E���f�(hѩќ��c �����;��$�p��Jܮ��{I�������fo�D���-8�7s�631� @u&�^ï���]� =	{��r��������ኰ���X����b�t�[�TG��p���ۉ����nT�9��,E��6�|���A��]O�ZI�U�O�612`���M�T���83wA�b���̾G�O�`^j��T�
t��\����(�;��3�)�x�=ӻ��Ȁ���*�����)q����q���d�����1�j/ͮ��eˀAY70*=秈����>dI�[�9�mus^�'�q�_~l\jl�a��X��;�����Ag�`v�L�1��wض�辤ꑍUe3�zQ��F��?ȗ�*�LM�V�?[�}��RX����,����>i�Kf,.`��@� H����i#���h��*Q����L����u'eh�r��3���;G  
��Cl`AؿqW/%d�'��(�S�����O'O_��V/zߌ[���ImJ��Vh��:�Z�07>���6�[�V4ͅ[�@t��?g�Bt��E�|�/��q����,���O��!ǀaІ(�*3#��׶�ʿ�:_̳�Mc��_BX�%��~���n)�7}d.���`�#�\b2�^}��.�UM;�*����0�җ�����\/c'��7y[���o��'RmVXʜl���`�&ȯ����F8꺛u�~��ш>�e�k��~�S���᪯�|}\��%�aֲ�+��a�l-l�Cf��vw\�������=D"��Og��"�����j���w�x��Nn��r}���N���F+Ж#�n�z��KO�9׽�kzY~�!RR�c:DAhV�MEE���~�\LMV᳆�W�ת��k�b�����K%�\���L~٢�
d�\q�6ptR~�UH��n��§�s��5&��B�r6I��k,�T�i�=r�g�'�|"���Q��%r�Z*�M*`��~����P��X��%$$W�8�Le�*�t�/�LR�톕J[.v��<xLa;��'AR��9�j�R_�9B!�ꛇ��"�JG�/>��W���2��}�M\��%Ƌ��|�%\��*`+�[����Z;��㖳�`��wT�R�<�nS�c���G���t3JQ�Om�Q���>�(��f��ݥ��)+� ^
����	�.)ۂ��!�8���v.�e�`0�����bٓ䍄R`�$�X4�|Ray�W�9I��O���<���mzw�ݣ�?�/��^ֹtO��26r��1�vK�=�<e�����H�
ŉ��i�+P���>�"��w��Jf���T�Yk8OY	�fQ?�%X��ɖc��2��tl�_���6[Y�#(�b#w��`_!���'R��Y1e� ���e��y�|4���<�ʕt�� /0�m+��0�\���c&t��ko��y�F�l2����\E�����WtI'Bْ Mڄ�\L��0r�lQ�l�^��-)�Pl�zJ�2�Gʕqʅ�K}4�	�� 6�5wC�[��e5�<$�8Y?��Z;���������0$~cd��&�")��ȰV�'�4��K/��{|)�:�N�H�۾NsM��X�\#o�'��"G��^�å-vJ��&'*�{VQ���g�
�$Y�sO��8��q���I�%�;G�*�#�v}H��)_��kZ=)�C��@(K����������q4�k�+�S/*y�0c65���[DK���3�s|W�q���\@��(�/lǱ�M��kVOMz��J
&dp?�<��N��ڪ��MP�6�ǭ��H�O)�٪Y��%�����@z"(���m�M2�Q�7�5)*�.�/�X�z{��~�O����)!��w{s?�h��!v�|���}�(�\X��eD�j�[�d6����+��O`X.VL�z����~h��Uhʉ�[чVi�x���!�B�4ݒ�	(��D�s�	��0|]N����v�M�.���{��j``�L��;�iY\v��jgxp}z�c4 ����	}�	*<TS�Z���#��~{�P4��U���� �>P��9]~�[��C���o�-K.ּ�V��a_��ֆ����!}9�/���t����ɇ�4�$���R�C}�`���*�mB����-���p^k�4u��&��O�Ͱq 1��_^u��JP�7O_������ɑN�����{�TY{�i��5^ܯKJ~�VB�s�?�A?�4"G>�́�2	�W�r���.�		=�n�o��:gy���@��FB2)��X,6���G��)�Ͷ�	4]V�u-p�ǉ8��#�m{��A(�%YQ�yl�*6����A &��
��O� �����J�a)d��2$2O���-U_/j�?]��VMf:58�x�2���H�H�r�H��^T�� a�Je��x	0GTS��Vr�y�p�y�$$�",_HC4�)cQ�*�z����P׌�~�����P���6�4A�����/����Y2<�S�LQ�P�w��m�|��a�O"�k�o�����[R�3�Z�?,�:�����<�^�ޖA�GR݉�V���4����1&"�;�\��_���4�i!��xG�Za���n֛��$d#S�K�������uhjnr�iz��n���ԠX�R}c	n4����y^>�b�Z)��9�+�-�פ��C��z'[�V�����R�] ���,�ʾ,3
 .��%"iU��n��
�;�/���w�[�?�%��ZU���>%�%�D��eI^�z�i���
��(���1�Pۮ�ƐT7���c��1ö��G�k���m��\(cxa۽�'M0�b�1�A��>��~� � ��@��&�Y��Ty��V������s�����Z~k�])���Mх�ܴ}q��8U:���uAc���lEwB�9ʳ�58!IǪ�'�xVQB5kv�֝|��l�M����`��q?;��B���`�:�DA�J0T�I����"Tj����-]��T���>G��]B^����8�kMJՖ�Բ�a�eb
w�@|��,\��4B�/79�	�Z(��U��C��T��جXN��S/h؆��J���ĕ��Ƥ)�H��~z��Ж,�� 	�z�ۗ�u��M�h|�s���B�TE�v�� ���c�
�h|i����z��}�V��1)����=o*[�"p{� �Pa
1�ow��T��=��P��,W;ɱ2y4	$\̘�T0E����^�T%Wn��`�$�����@�깼ٽ uu�<=B���]G���b-ZTԠ���9ׂ�A�Y,8[k�=ֈ��� �aY�|�9
e�aR80���.m8N�� <̫��ǖ�9��2�R{���s624���.�*S5 ���֯s��)���B{�L��`Y�p*љ(|���@]��꒮��կ�l3���U�����R�^^�^����9�;�_ȩ7Jڻ�'�|gXL�V�< �W'~�ba9V��PU�7Y��,�t(���s��Ӌ�;P �����d�-"�h`�>�A[���D���W��l��';2�M#+��zțc��s9=� U=���C&z��<��T��T�CI?��w���,��3�R2�@/0��ߩ�u��rfW�+k���Y��^hiC����gl|�N֫qz�8�Ԙ��� �Ƙ���fARq��nPLS�]ט�\��n����s���X�Y�E��17������j�Q�C���h����NX���h'Q�%�;h���BT�ۈCH�z�hݮz�=��'<0;�d]��F�F\��Xu D�X�\tm����)kQ��[�[~��<�!��oɈ�L끼���~�9����Eޣv�6�1����}������ۖ�����b����kuՋ��L��!]���r��z��T^���탩�#k�e?��HFJA�	�	RQ���Q��F���Ab�)�(Ț-A��Y����X�+�Ź�_�3�s�~��B b�X��6��%�j��-����DE����L�Jx2�#�{�#�p���<ʭ А���ˣ�X�U�VΠ�]Q�G��.;�U��u�E����1g�L��ٖ�_�������a0m�xQ�S�F�-^Ƙ<��q��4�s�l�]j�r�h��$g��v��\;�p��z����鑧QZXe�@�p�IR�9qZ���m�)I����lH��c�I�ڂܶ�D�0���1٠�Y����p�~�u�I+��'�%xu��^�}�X��E��+��j�v����J,��8c��r���[{-bd`�܌��X*�:Bn(?�����#9�S�@�Z}I;n����x.1��h%+hng�ϳv��RQw@d��xZo9�[�_�8�0|���fa`=�qr�~K�( ����{�?W��mÚ�'Idx`V�g�������U����m��������O=N�cðT<�����.E�'�Ɂf'{5��M�D+kBD��3�߫�U����<NF4�)<�+�.�8��pne���L�!��/:C����t����O�Y��"�A@��T�ŃMU������ֶ|��:̮��. ���$����L���t{����07�o�$"�c���>��m��4g�u��S�F'�o��K���vY��>����J_*�(�`�y���3�j��j����n^�G����u&��V���R"�5RR��+ !d_ɜe���zջq��P�S��� $�΄x��S���VԊ��a-�P���Qc��������'^���/'Z����On�$}��5'���;S~K���b�iNE��X��&A�?�^�L%�s�ƕ��N�!��	��$m�,�3H���/3�|�][i�d����`�����Ž�?ҁy9E���ȕ��VI�YH)�H3�% s�>�������ƉF��Ч+�\rG'k.7����SCfβ �y70�>
֊g�K¨�X��n�̈́��T�{6��K)߼�-�������@�(=�F�̍��E�����roQeUԇ<��y���.2�X��ϘP��"�_f�/#�v���;��n����Čsp��k�H��e|?}��픓�"%���\�M㨸��>���9DR0��d*ى��a�n��*Io������|�WP�^3���)�\����ulylz�R*a��Ʃf�*��b��t}]�Y[b�h̫G1���e���Q�7��\<m�'Ȳ�F��$��E�'�b�mc�����}��N���l�]zD=�1qmM�m�`ܘ�2;��OI�����$� �(A8��~es�e�9)�x��U�P<�1%Ln�X���Ӊy ��Iw��%q��\rKD��xZ�p2_QC����ĝ�LVY�u��#�f0P}���^9,Q�\O��T�^�p//��]h������xA�y�f0Y������	��G5t_�ƈ�]+Ԓ5��
�+oN�-�:=�Cg��|O��>jkE��($��^�MC�ңyt�ŮD����w��d\ĸ�:&��<ҧ�M�ћ��R�&
���s �xʒj0yY�nx�?�&��(�=�nz^����2��Ϣ
Z��p��&+�ݰ\�NǠ�`�l�~F��%L���mO~j<��`���f���:�Ԁt��� ,�x�B�VI�г��k��CT�L'�M�q���kev�i�0�O3:��eИ��ffB����P�W�ڢLE�X��LuԱt��f���b�/n�yS������"�N���݉v�R>M��sT��t����cl_P*2Y��x�f���b��Iݳ�8>��J����?J�}j7XJ�טN���\<�UF/�*6�ǈҬ�KU�vr��%:1#��x9rE�D������F1�����nΎ���Bj
n�Z�O��h�2���DlLn�A�<LwAh3�D:��Af�	�%8c���9����1��M�BL���&���CS���ٱ�����t��K�Ŕn  m�� ~�R��=G[<k��y=D+I�nTu��5IPd8�*���_����4s� �+? D�le�����05�����^����59azc�嬧�K՛_�|�������I�E/�8��<έ4���Į1>�:�
��Q����]���t�v�|i\(L)�4m��`rj�m��UW�>D(b�_������R�(ft��;!V]��T8@�΂H�b�fJІO)�@뵊Eg��7tD��?���&|�P5�>�dG*�h'� ζ�tk����F��V��ER���!�<�J��Mp�ڟ���T-���}ش����f�8슅<��z��a�ݙ�1j�d�Gk*�z���{x@����41��P:O�^Q�8��M���24�t(���.��S�Mn��S�z[Jxٞj�NB��Y{D�ZzRp�"�F�����8�Loe��:y��,P�5�i{��w4.N���o�DG�P+g�V��al��m�xA�{�w�a��=�}>��f:�^�'ંT��6׳F�γ��&����q�q4u��!��/�\=�ҫ�QZ�+e'� -�[�A�����JCp�7p��E�&-D��7��X���+�y����ai�m���_���iW7e���ӣ��#k���*���j��ǃ�8���6ՔKA�RWqv��I�n��O���}{>�PSM���i��6
7m��Ћ�\/�oWԑ����#���2liƅ�tpU���4�~�;^��l�p�	.ތ�zM�(�G��E�R�=�9!��k[3�T�5g��iR�h k{��gh3���6��Uę�Ř;�ʆ9�3O�"�`8`�ϖ�C�0��L4ˮ
�+)���J��/[�6��s������@�*���]��I����b� CW����O�:�@d��\K��+*"�I_��J~~�͑�4��n��Dc�A����ս0����ߺ�$H�Pe�eVi~%�{�)BP<z��ĝ�x� N)jb�u3,<
xF����^��9�B�+碞*N_^����²�6����ޗ��]�����P&�K"H�F*13��~|��]���Ȣ��f���||*[W��tlѓ�|����ۘ���c 	�L��u�f�g��n��;�MBlzg+�k\�u��KO�u�,�9�>�R.���:{e�����  wr�>'"�L��<Q�x�eI�R����ν�i#4͐E� ��8��'�J���5����3�9����h�� �?���;l+��D�z\���x%5�c��D�̸�]�8OjA,�6�C��+�S�����Jt�FaY:��M�N��Rih�4A����I�k�>M�K_6��� lp�4��3�)]|B���l�u;��ԧ9Θ���dЙ��1�z=۞9ƿ�X��m�~a`���Ǥ��n�S >߇��:��Z�?�aͱ}A�q a�)�g���Z@�%H��sQ�c��5�A(]��s]����"�Ǫ�q�&���XYjX�$w>���/8����&��X)�p�go�.#BX��Qu��p��)�3�#� �%�0uJ��m��m*.�o@��A�ۺ6���6�$�7Oz.מ�])�p�_��ps$i�֯��^Gt�f��&A�"ܰ4*�$]��=��8�/����h�q�z�4�*���2,	j�ʑ����[�i� ���������&O��<��}H����B�K��ã�+�N�OޱN�{����E�L�|Y�x�Rx`Cq�;nDe��
ŭ=gh�9����muI)-TU$��u��4A�Y�Ѥ�{@Rͧ`S��(�h��p�˻�����G?��[ Sj�_N���2g���\k�!�;�BN[���{�t�(p�tƗ����#�ܒ<|/���zv%�ȥ��ٗ2�ޑM���書��;8������m}�poJ��!�F:�4�-�!���&2Y�������&�Q���LR}�
<ӎ˾�I��v,U�X�[�N^�i:*%��7�5+�EQ��;�{C��(? �}��&�A��ν�`t���9ޯ����o����Q��L�{S���L��&Ƣ��������t��SB��X,-8.Egz�y�	������ד�{KbYF8��!k��#:�/d���c4�t>�5������{d��E�������B#��V��y?��=)�T?�[�Ă�w�� �`^e�.d}|�=(��?�y��F*���kp�ٯ�y�B�X����os\���Vy��� |7����$�֥�2�a|��E��l�su
i���jV�P�b�W���PkM(�����#Z�ӄ,rT�c9��y��q�3�K�-|E�V�l�qIT��	E2�y�~��qg]�A�xc��>?����<o&a����5ao+įi����`���i{�Z�B���6RRP�p;���*���f��Gݔ��c�\�����`e��S�Ɓ��y(L %(g?���GjFmYv�c�[P8��*��Enb�lþ�Ҕ_�g��w}�Gn�ǜ����-x?=�DgI�I�T�S�F4i��^|��7���7�����kch�'����$��_2����I�pk���P�͍��)q��7��-YC��͉�Úƫ��e7�%jA��->,,>�J��ohp�O�@+��D��G콡=�ޒ�<a�p��̥X19�9ۡ^le_6a�{-H�~������bJ-��Ԥ�]^����4̤O�1�9���T�����q/��5VwH�(~�i���Q0д�bV,�y�ھ�r����ʁN�#&f)8�(�ǃ#���^��5VpC+u�`�D�����go�v�-!�8��=���Б�����v)�l��
��Ahg�_�9�t�7{Gb�#fP�1{��v�����5�+�=���ȉt}5eZ@�ߋ���_�}�˝"OJx�
 ig���â�2Yx���R��PG�������d����Xۃ"��ȴ��.�ֹ��ܫԗ"��m��3I�3�*�
[��ѿk>h�=��>�� �����[G���3ۓ���oJ%W�&�)�8F����9��m�b�d��Q:t=�(�4����h�f%����Q[]�?�=�h�N_�K�>΂خ���W�I�M�c�����~r��lbD�E �J�af}�QT1@�N������<���TE�\q*�-�b�C�1�($[���ݴ���1��p��xx�u����`�_Ǻ�R����+'XY�Y��m�'�q�2�	���jpQ�����e�
ty��Gᢿ5z�M�P�v0)�K`�����
���k7����E�-�"Xr��5��G�_s]3§'G@��m+3}j?�=�?��Z�9�D5:�HH���7�|��@2�(���C��(_�e�ҩ^�hu��֩���:a�(͕�~2��[*��[8k?�?,�� ��xmb����s
Pr��5v��y��'	~<	��X�eE*,���U�r4�R�NHD ���9i�=b/9�$���~�d9ȖR�x+�C��q]�������rE��^&�%em����j���̰3��b%����bb�v�x��do�m�E��>��N9��O?j��|�4�؜�+�3ۈ^/����L-�܄�.��!��Y�`F�}5���*7^��Bo�ng�,�"���y��-EeyLf�A��ǹZu(�2C1*��|瑮���+���.CP�#��=>��߬����wh�'��f� ��`�0�x��t;�Mg.���������K�%E\T��N�
7"�J���5��.�hF$�%�k�P�/�>���{���O}A�Q��O��q+�þ�8w��q i����u�\՝��p�۾�2���h|�o�����1����@x��X1c�
�E�����g]�ށ�����%����c���Tڶp ϔ�nj8�N݈�������	��y?�#f�1i/@2�C��1�ֽ$Wd�$�������o�:���aI����0=a�M���q��R�eu�r9�Q�c��(��
��{�ߢZ�!��Gg.��O�'�c$y����^N*�loe���W���6F�,�z�0kr�	��o��K�B��(�KP�l5r��&t�q:�_ɋg|�tKq���	�/Ň�E� �h����]��#��r	v0����2�{��B��E���l^ �W�m�N]��ކY��ᬭ8�tkO�Ғ��\����C�����Al@���HLK��&G{�&�6��n��^�޷1�����s�sMe��6v�Fr��I�I���$���/�"����c�2�ͼ���o��aud�8��*��������1�r~�Cn������&qk���r�2�����(�7��d/�� �,�-1ZU<Al��K�u�J�tsO�̻�[a���ӓe���)8S|ԑ�4r����a���	;00"���	�IcQ_��,n��P^���s�Sʽ�^ʸ��z�E�[替b�������{{�U�v�G�n��, fu��Ȁ�9���t`j��*���y�gt\�5>3����2�{��O�H�n�Ҿ<����W�g��s,2�=$��u�g�$�AJ�']�-���@'��(��7c8oz�ށcv��,�ʮ�\]�L��`Q�`��)����р�X���2KH�Se��GEo;6����y�U��AS��v���{�:���n�	b�,>qDǳB����1�;��Z�4�E,\��h
��~��]i;,-��vL�A�f��G��&�j�Eĉe	X�q?M=��,��0y5+	��33�;�]̵{�_'@|R�}�1���ٷp��!�-)��('��#p�t�v�÷�xo����u����*�hwY�=R�K�}70�+��C��"z�]輓�ui���RGaK��#(���D�� �
�!�$7�d�J�L�lo� ���o`Ύ)��i#i-6��,��Z�x�JqN"�/�Cx�FgwR3;�8�Nw�� �E�N��T�pX��,w�[|,�Pw�LW�������xvip';�������3��&o�y��;�NO�/��+[�^#M �"�5pq���I��~$�� S����H�*4x�{)K�����Y�@Ħ'Dk�Nk~�I	y���2�rh-[��O*U���GM.�XCsI��P�BQI�aQ�'{�L
��X����<�tS��_�Ӣ��P��w?�F�2p~�T� vI� N��~h�s�;e`���
�H&t����5��u�4FO=�J�2�H	�t9�Y>deʨh���|�)D�A#k˫��ϑ��y$"޲%&&*T!$��L�g��@⋰�8�$��
+p�0b��~ix2���⺃��E�ǟ`A�E��F5dt��%�cf���ԋV㖬C�g1Ʋ�(�ݼ��"�u�Ǆ�Mi�h c#l0�fcq�lx��.�Zg�ǖK���'x���pݱ��)OT0-:����69��;��*�A4B�� �t���x �]�W�?����;���|zA���(g۪�!/��nX 	������*p����o���|������tn�+4�(D���p9���3˶��I'�bBτ�Sк%�F���m�A��:2бG��k��N-�I���]�:z*����d������y���|j�k/�%L*ו+��1� ���o?jজ�ΫzS�����=�݅�ZT����֌=����=�D\J���+�����9��K��M�+tݱ�?��y��eڤ��F�Q-���Iztl50� mt��QG��N��#Y�Bnn;S+ޭg��}�FS�b�$K���ЕW	G�Gj�^��)���w�; 鐈�)=*N���@��V#U�6T/i��rT�3�f���~$��u4:��0o�f�%P�� � �����걄�l�(�V��xe2�S�� ��u`�%��~�a��%�]� p�!vμ6����{��
��R��*^�k4�h�BF26�.W�c�3¶r���(�!-�+q �]}T@xsB�;��n����h6���`M����v,'���tsJ���1C���Jܷ�v��gŒ��e����������.9�6O�����8̦�m���TQ#����a� �,m���0���:�Ȝ�����&jP§�1��魊W�踕�� �����b���4]f:��2e/����2mu��������X%��9�hT�)�zd��ɝ��;�佪��1�L��|e&��E}�eN��
��?���Ƭ�>���	m|�����-9K��-|<Zy��C��� ��B%��w��3�Ν.�F{p���'#Bz�Uw
x�LE�̙��r�#3�:��$5�@z%v���`P�z��b����يM�A�B�~��1��I^6ZD��<�`�*�a�W�:߫��~>}���{i�_��S�Ը�;�I?�~=�������̐�$��a�?t���6_7sGy�!yERR�:St�<@p	�"֑�FW9B� ����_�j$ͩuW�7d/��L�=c.K��|Ag�w����7JO�� e��i�S�Hc�i�<j�����5�������8G������@��~"9۰�b)hm��l�ҫo!i��L�phg��U-_(&� n��ʼ����#��#'��2b��
��I�E缺�}gS]��Z뢴5z%����>9%@5��F"MUĭ]���a�-�M�����f_��z}�q3OS�ҙ�V���i/3X[ �)y�	ֵ���5�(ԧg:�o.\cL1M^m��xA��k��`Ux��,j���+|п��{e�2�Yx@��b�ѵ�	�DB�Z�����QCi��CD��Y�V��	Bʂ�#j۷�G|���K�5ǅ
 	�j��B��\�*�,�/2�x;9����vޛl�hv��������iKQ^�	-nE�>�O�w��]B[{�j���:��)��9��[��"Ƒ�RS�k�ݦd&"��z����Q~�/:����A��?��:t����ʘ�B.%���b���B�9���ӏay��5�6?��N� f������i-(�{�/�7QC,�s;	G��26��Z��V_X���0șD�cV$��#mf���S�c��ˡU��,ȿ������wǳ"�5������\tz~	!fz�¥���`�cP]Z�+����=��T��$�J�T�� S�܅�fK}�(��C���E^��P�'�
�GX�؀�'��D�1�r?@�`*���`��I��N��
�x����*�<'��Y�Q���8�u���88�*j=���X�i�ށ9�@gJ�<��>7$%�&�-�k��ot�6��kŇ8�8��S��EӞ1N3�#���@��a
���7p�V��:3��2��� o�k/���,bYfY��S���}�\D��F��%�!4�M�\�yT�E�Q��K��������T,]b�Z���ҝJs?�;5�Xn|h�B���WS��I� �R,
�$g�KܢT�8벝����鎁lh��&c�{)r���1��ȟ�?%�2Z�:�)��꿘UH� �x��w�;fی�rȊ��-�}���L�մ�C5�*���������:,Lv\���+ZQ��P4� *�sNl5:�����3����?q�E�z�.�~č$RMU�q�4��I�ڣ��J�ک	[��e��=��G�<b�o�)�{=���ԻB��Ɲi���cB>�R]����$�%�Z!3$���\�dXO֠�$�b.q�B��g*�Qw�Pˀ˚��3�.i�uu���ޭo�|���HV:��Li1�4�D��e��\������f��3�D4�����M���� r答 4%h�KxV�����QE��b���}��P��X.��G�  '�{�M�Uv�(��T}2-B�Ѩyf�B�ky�k��V ��.�Q�Fi�G%��X~��@�䆜��SQ(,����{��������Ǆ�2�*��{;s��3#�8)Z�J�$��������<���n��O*����c��d��S5\czsT��F�w<�C�T�������1*��g۵�g)�n�2�[�`��_v��[�CH���Y��X�0����3���Xh���lJy��7$��;����'��7¢F�b�غj��v���r\�4�O�9�J[K�١yРvO���C��B��&[�K��t�lM_(bh�t�YD,}����*��Xђ`4*�}�㸼�2���u���N���l8M���r��d�����ˈ���B ������l;%1�0�2�M�廋E)����3	HB̲�#�5-fnw�&�OȍXE1i�_�T��V,5�����G��>#`fǛ���D�w�luY�!�!v�p`�>��G�$	�؎:r	)��Et����@\P�o���������8�)\���ƭ����jh�~B:3���ۉ��M%�h]��`H�$
	���e+�i����)�p��8�����;P��4XY���ZG�&�2����9��/�6m�o�-�!<�[��v��~��%�ک�ܫ��K*E��-�6|U�7��4]��P����UB]G'h�8b���/=���x�j�E-d�u���#���~3?�q�%��m�x	^
.;3ѝ����0����Zu�H�6XKlGv�}̕v4Cp�7�n���T�Ʈ���z�S���٦ T8i�)w}˗�ɮ"�~�z�&�Y��f��;��Fc$عɮcF��E�L���~V8�_c�;�)o�m2�l/�s�{~���vkP����Q��OI6V��m����õ.��7(r��=�W�u�L:s� ��R0s�M�Y��.��B8�Z�.BnČ`�x��m��t�;xtkq��.R($���@$f(�@+�p�;?��������<5k�36TU�;�AЮ+*"?��=ډx���	�~��.�-����K�'�`s���ο������`�;œu�vH��~�%��?�1�SF���v�2�zЎ�}�u^I���o���c>�/c���?��T���RE�����B-��.О�n��緵D$����G5J��cC);C�N��s0u��#C/�$���e�ƌ��>��ߛQb���0�-��r����\�!I���S�G'mRX�2�yE�[�K��'�k��z^����y��-�$EVD�˫HKKz�z��j�"F���*�PL����S� < Z3��_����;;�[}dcr
!�e~�N�;Tu��d��^_2\���kIS��Jw0���tv�����&�� 5]" �~����k=������2��#���@��P�jh����3�
f��Q.=�s����š8��cK��x]�{����P�!&�wj% P�^��9�N�Q������0���bI��	^��dM��p��V�4ɝr!�xֱ�xg6��Rm��`x��E�3cr�G�������S���"�U����k�U. OX�׻N��lu�z#\(x��\�˲n�T�"��F�ؔ�}*��	u�Hc#��p�U*�� ��-H���dS�e	�`��� s�����ƭ����'�Z2�v�e�S�F��l%Gy���/��߱��]�-o[x9?�k�߇U�]X��ߒPQ���¢A���zhm�#3���><�)��q���l8����+�.�K��H�%�9�{#�JY���@�^����z�\�;q�l�fB�O�n��>gO3�l|���F��1����C�He���n�@�#l��a1q��t��΃��N�Ih0�>A��$s��o
w��xPu�8��:�T,%x�E�i7�����[x��p��dQ҈�@�7���t�n�k�Ō$�W�}%&=�,D`��@��p&K�� �u�P�Fl��<L��$�8�ʓ��Z�^�X4X*Pɳ�2d��ބ]^�\��뼔'>?�\�h@Aq��2����ȵE��IC!W�b�[:�͓)�F�i��yTY '-L�/
��:�z��H��!(
�p #�����~3|�#���d
��55��(�B�}��\��A2�v҄���W{�8�*�ff��
�b6 �.���o���r6ϑ'/z�|�ؼ��^?/.���a��QˇrtA������	�93�=�m�J���s�-��C���4���k����G�-F'�/��I���N��|O(�V`}[���/|�KR~�M+�␋�su&��5�u%��9(�hl&���K\.�kgk��nSw(?w-P�!x!><�L@r=}&�K��V�,+���9԰1	xf�s	y$��	�D�M�2��S�R��Gt/EG���M**� �q�f�t��/\�	�1�E�6fϸ=���q����Ybd��۷v� ���{4�Mlf}U���I&�}�U%A��=�P_�G�_���erI��&69˧ �P��G6��^r���r��E�6��]�%O��6��V����؀�vߩo�s��>L!�z`�Hܽ~0��Ji�����p&y"1��MXBX�n�%�!��&��?_tΠ~E��-܄��(%�e�
��
�Iq��R�h�}�]cA�ɲ�\I^��q	�T�.L�����*ă"�,��n~��k*G��F[{��0ia�.i�⟉"|UuS��C���o�����L�Dm���i&�o@n��f�&8���� ͽ��JQ�!6'����Z�����Z����|��Wb=��������
P�$�K���s�@�ù/�C��0���^@�˞'�;T��R����֔	u�"�K9:�ɹxz4����(�H�u��"��JXW�=������D�M޺��_�)A=�4J�#��m�O %?s������܎J���]!�H��na�·�f����1n��/R|��/�mg��V��P�����Q�m��u��ݩ���x�9� a�p�e��H�ZH�|;ł< ����ۧ$\�RI>]S$Dd2��g<Zw&�o��bm�ͷ�%^q�f��ў[Q���,"��<tz�����m�&��pTL��g��B���Uw`Ϯ	����a���NE����T#�(��2�4�%�,"��3�.w�W<N� ��2�r�=��h��t
��o
���SL��Y8�ס�������S
���20�YJDAb���8��,�+-��bG�;8�s��T	����Ă�Ѷ%B����P�*���A�3^)b�8�D��_mV�=�][4���ms�������_���K�y����)�Ք��&���e�p������1ү�w��r��{W<77�K#?�10��;d����m��r��+���[���5<%uau��SLz���R�lZ�+���T.{�{��^�0"#�	Y\�'X"�l�V�	�o�]�X{��������`�@խ��*4l�nO���SI�E���6<��m�?Ou��n6e_��0t�����QS��Vu.�'�TЪd��ۇl��`��7õǍ8�\����J���E��| Y`�уs�m<	��d���c����y�@��Ѿ������@�0:]�P�J0�Rx��bW'I�30����_8O���{Ԡ�vRsB�ם�q�l�|�w=a��S�;Kx׀�8<��2��L>��_��q@Cm�cQw�Q����1�3j9Dʋ$��d��:�
���Ѧ����h������Ø�z�T_x�����%�-&b�IG����g2S�Eƾ���}d��Y_��։Qp��{%���¤Ns
a�J ��a���GϽ����K�Ҏ��O��@W����Iǈ�:ݓ��ko�`~Z�d
����@j�~V�9Č��b��
�D$��$������
!����������*뷪e7�[��5�o?x��������F�(K����������P>tI�@ɀ���L��	I�"�h����o��p��Y8@��g�	�!���mB��Fo��6'ER�;��~��K�<<j����Pa�PA����}�m��t�ְ���|8�d�hڴ.iJJׁd����6�:����z���-_����%%�}���β%��h�]nc,���|���'�
�!�"~��W��3�w��d�J|�@��C�N�<� ��9����M���$;� ���}X�+GHB����PrqA�H�?*����v*B�_J����93W|pf�"_�i��A�w�c6�1���b�B�Z����<J�8c�(Z� s��DUS8f�<����r�hH�	�\�4��q<�ג6R�B��–�!M�:�J�1��|O�{��ՆIc5��O8����2����9�7&g;4wNi��a[o �D��0RhYv�2���)��6:8��e:�f����1�2i)L�V�1<@���˱4b�ܖښ-L��9�-�a��։�%�%&��g���||)�~j�W��G�s����N�=n�,!k �{̓��Js��g:݀�joy�ɘ�d ����Z^�xb�B�<1�0q %Q�L2��t��mc����	�5��/u<��֡����z��4�7�5T��whLV��y`h�~UP�e�Ѥ#s>}��!�T�32�)[��SY�.�t��t�|�N��b�l��p|_?<J�e*�C'�,�uy��~+�L��~���믌&���CѴA���v��`AA|�6����:P���/}����
�`Ga�c`^�`wU�Ww&f.�U١\wl��B�~PX5V�Ir��d�u��/�-f�,J_ʏ�� �}5�+[u�n���8��h^��tߏ�S���r}� 1�Z]�	�g(�Z�^�%�4��xi�xф�9���0KN|`��~h�S�ᘥ�4���� y��{���@#J��󩋷�]%:��C�}i8�yU�(��$��y��}��=��'��u�[m���cG�,g����)�`��O?L.?)����Kt�x>��f�ψ��$hx�e�s��[�3L�6i#�!MWxW�;v2��Ok@��aY�K}3��T~��[C~��a��t*��׎�*=����ZX�t��(�I/�w��;v1V�A���1셖"�Wū��-6;Ab[��i$j��?��Q���I���x-a�/�z��6"R'] ���p��49������+��:��G���jG"�nH]��s/������%���qO-(Z�1�	���ߍ<�p���������j�� D�����۶�a��}��Pc�@�~�6���Ekk�)�h�eY�W&�J:���'�5%�]8�&�R��'g_;RP;�����&�+���:7D_Z��hJB"1N�<Y��FŘxE�Mr�ْ�G����<B#���Y4�e��]�[1x���#(��Ƃ*��5��]�:��9P�}���zZ�j�v�'�l N��{D��W��(�@+�7��j��&2�0�p�گ{ӝ�� |��zڣ�ZH��ZP�\�;�=�(��,E�pF���t���m.Kt2n���*���z�U��ݯ�p������=��yf�r2���o��]��&������T��P<F!*̵㏪A�\�"���F��ǩ
�:"�L��_lۄ�qA�6������������*���>U1�rg-�~����3����q��l�ȢG�k]��(U�c��E��X��������}�����@7`����0M�nG�ɬ]��.�������Ÿ�s!��ԫ@N-ܬ��8�u�;����)Q��(L�.�h�������3��v�P��x���v�V!Ӓ��g?���@(WG+K�V����_�y=4WJ���5m&��WNy#dD�J:v<�>&A���h�F������~*�
�(#F+�������
�l�,��R\H�*�v�^�׎>��UЕAk����r�MbT@v����b�ƍ����jп��$�
�����`����}�)I~dQ�l�8�J!��|��u7��.]F�,���*6�^@��ӽ�+p�L�c�2EЁ�L�1���5j:i(+�[��x��_!R;�r�BC��U�x�P����!��r!�L�p=��q���ێ{ƴ �ɴ�����ؕx��Y6�}UaP�_	��V�2H2cqta�yP.,��?�	d�H,����%/��2�[���g��^�m����ʫ�eGS��Ù ��+1�Nŵ#��@Q�>�^����'��8�K6 [�¼i�k��`>m`�� 8@~D��#hf�����E	H��٪��1�|�x|E�Z�8k�l]1-���i& X����l��&hj�����TI�|>�I�b�J���Qg�ޮ^��O����P��g���n���dh9��0��m�ο�~�0xf?ت/�yݦ�'���vz�R�������c{���{atS�̼���xh��㫀wayˮ/��< �oҒ'k����ì��2wY|�wl����r�rwW���捫�f�-W�;gM�-W��,����ϭ�z�qc�\�|���Q�-�\��#���S6��[���ĭ4�q�I�{��c�Z�ZR��*�h�����<9�j.�j:O�eϘyŉKN�=.���5���?�jl�:i�Ѻ��|h_9�����b�.�&a��#A;\��n�q������wbqa�t��ٗ��)���=���g7�>d��7��/Ю.���`�5�E�k�ש?d<�<�-�p�;x��J���C=�?&�!���*w�b@l��c� ��(�J)D��9H��=^q������p�_HpH���d����	��xFk\�t�<Oئbޣ�t_����f���-�O���iL]Ѿ�:�T�� >���:�Fne7A,��:�+����&����Y���7��&���I{W)�/PD��|�0d9������#>��h�	��<Q�dΕ�g��\ ת�*ț<~/K�R����Мx'��}��}����Bvd�] �/�Ț��(��)��Aɻ_��������)�n�J=�th�D��N���6P�$�W\vC:Zܡ��!T������d]��o�N!�+��0Þ0�PU�i��L��u<_�t��c��!&^�4��E�K�ݒ����D3�e�����3QRB��g�{�L;"�'D\���]��t���^�0�j���.y���=9
Wc+��4_���Ѳ���3�j��y��Ƃ�����&��Sk3�m���u��w����� ��~y>���tk�ʞ�rd�+E�j�$m���y��O���Q��w����!�j��q��zD��X#��FB z�C�Hqݐ�܏���~]Oy�2MF�i�B���+��NqWJYԉ��-����(�M��E(�PｅnYB��>��� �����c��"���#(oo�RԲ^Ff,���6F����èh[),�F:�{3�j���w>���%�S���?�[Q[�N>�쯝�̻�m��9( ���!҇&�O*yiN�����-�|�x��o�>�9KxX�HG?��/�]KId� ���kY��	���|̡�������rk?ͦTr�
-]s�z�S��T�E�h�	?ň�y��~]\���W�<���eXc�#��������bȑ��%5?q�]��^Tң��B�{���$�q�p�u���$�g���w����G����F��)e6��;�w��xp&bÄ�n��t��8P�7�w��DNe{��,>�QTH�ƆGɧ�1�FFD|4̟����`w9<]
�6>���UVU!�#�|�&9����!�@��a��%��q�"�Z+\LaID�,��*z��< ����
e8��pT��1��/܀*u�w�#K�@$X۰ץB+2���:r�!�Gjx�7kVx/Q�Q���0Oj�×-rc�D"�����&Pk����)� F��,jeP�X��5�o8Sl��a��hd�D�O�ǌ}��c�Ж;��v����:'�GZ���z�ד<eci������oQ�9�`̐%�®F�+�#�]�A����vh�C���D�]x���H�RǴZ0� h �y�j\׽H��w��B��>K�X��S����|�k�/��&�T����k'κ=T���� %j~������IIP��28-�P��yɫ�D��7�J��gF�p�pu����%����B���ۯ1�Q.����~�}�*]�e�1� �z\N�S���Ƶ�/������P�~K��(��oϏ�$z�)ٮM`��zZ��_�[�F��RQ����o�9Ip��f#�6���7�3�J��NY�;���a�Tx�+~a1��.��>��&���^�hD�$9?�	T81@�7?��0�-��8��Mr��b+N���`(ZN����>�ٵfp՛"�w$ o�����r(F�zH�|8�Q�l��I��n�"�:N�e3��_ �$pYK\�Sjs�ʓ�s;�$,�-�G��?P1�?(Er��������H6eQ�܈5�ү���Q�F��#�X� ��E���%
ɧ����-�^����3[���]Uw���P���L�z3���D"Ҵ��n�S4��ϭ�S�P�Ϻ���K��;Կ=��_�{y���b�@Y��Q�<ÒT�X���Dc��t��������A��O�kNtN��x 5�^��ѷ�_@$��L,�w8� &(<���2mec�NVe���k��5�8Y���R��t��.aX����,u�>�u�:ޓz>�B,��AFŧ��;�jw�G�Z����J�S�?�u	�ӊLf�Gy�~*I]��g��x2B��U�d�� 5���w���c2�#���S�����DZ#�Σ�s�c_�M�D����ɛe6h�5��}H����y0^�XV��!�a�y�v1�͸�,�csk:}���I <�/�'1\��ܧ�d����][4q C����M��5�����(GߛGE$�5Ƣ��*�H`��{�O����Db�P�)��6���)�`SO_��k�cA+w@��e��o4�eƀ`#g���w�&w�b|���j�eyy�uP<[���[�x���<ܢX����jA�)$�`�cj�ĠC̜�RWv(����l<$4�6/'?�W$0u�QkM�h��v�:�
��K��C���ɶlc]3�����6�wE�7��y5J�d�vvD��P�[�y�����e��ب�%��#Î��	���٤��CM���>¨ka�y�j!>!�V������Yb&�H�D��LEB���E��\ Hx����.���� �H��O	��lU�W �XF�D,:�KX9�z��0{}_�`�7[#��U����D,�������c����R��8�F���OE�L�A@�\�o�΅�%:��1H-	��:����N�Q3}����8g�#�c���K��FA�������͊��0Q�$�0��-|���!k]����g�%�r�)��N\\�+lck�AW^�����Q����I�yۮ�[c��H����;Lf�J]d��>��тqD�\ �w�
�˵_���P>p�����(f3K����|�,�P�Γ���x=l����
�H��O�ʎ����BG���&ꞥ�m�ò��:�����Iv����*�-�`�A���.����{-u�O@(�{H�0�[��X���k�3'M�(�4;v]�0�E�ED3�L��*>
8�;��7s�!ѷ���[��vT��ე���۷�j�|�mh��3:$X$�����(�*D�dܡ)^��@��P¡)���1�`�L�w $R乂1k=�������lk��jm��<�0p!�q?�~nM�j��\�g�d����� ��~��u��|���������Iԏ��͈����$���4��p~����6.\^.��U�r\��A"En+\0����hn	M���A���Y�q�i_^��qR4}ɘȳ��{6�H�E65�_S��jBB�WP�I����Br3�U戍<:�J��Ud������!o�֚�����e�]�)F�(8�-(|�9w���(�L�`�'��5������M�Ic"!�Sdr���Q�rW��b�ht��E�3�z�X����:좊W�g��,g.�?4A��3��%��X)��'�;��%F���V}��"
��"�M�����Hݹi\9c=��"����\�1���دODr���\��C��ŗ����|���R���׉a�Dz>;��W�]��?{�ӈz1����V��o�Ę�8Z�����b����i,$<��g�i4h�!k��4.֝G��`@	n���R���:	U�H�23b��$�E�c{ �I�
�=?��ڃ���Ǡ�)yRV�]z�����`_gR�����������)3�����9�D�$ڸ����҆+�e������B����#�J�"R,@A��.s��]��*<s]�d~�����3|gL)��{PE�K��^��?w�t����^�Y�̌<^w`k֫b+G(��N\�%ZK_۸�����& �b?��U,�/髑$U�a2����K��:1-Q$,��A1�4�#���%�#��7���4<�O�ս��k��'R��Wv\k1ۙ�N)���NZ�7鬐!���#�=���7���@���&̙&_�`�]IO��9N����Aԍ�)W�>�&JP�B�B?�
������j�Pg�fƧ�1 �V�V��G���xD�;��-��׳�Wm��|�32ZОz�K���؅��(�3��1�����,��↝y/�~[Q��N��:G������/����g�zdN+�o�@~e%�C19L��q��7%�'�.h��+lp�Zffa�]tm�]2@w6Frܭ����a2]A>]��r�#�m��Y�x����WR��I���t@�I�m3h�נ]�t6�o�LZv��d<���ߜ�.�~U�)ʩ�ڗ����3| b�&)��L@bȕE�0v�◘+n�5v3�^y|>19�
^�!��@����s		����Q^*�b����@傳A��M�$���%����;�`<g�\��D�1y�fb!t%��%D�F���"ZOL&�^CU����F��W��BP�N �E��"��ꂱ`���|ՠ�=�sՠ����ҿ�メQ��f�a/��ZY�%���֐	[�N�����e�<��ƶ��$HyTg"A��J8�m�3�ԩB�6�\C��8:k�AA���q�:Q���+j�B"�r��N��4`���3^N����N�>�;e+�cØH��@�[�����-^�F6"p�����6��;�ܯ�_��"3-�֑!��Dx�P|�5��^jx`o�ʄ�8X9*\��G�[&�t6|X�i�v����E����E�I�%�#i,W%Mq��u���C����7�.�|��#�_s�v^�V�D�ޗ��4~�����4d��<�)xm�츫�O^=�3[���,l򥪛�2���nBI~R����rZ}���Ⱥ2�{ٚjDͤrw͙�
]�B���Ou��"�h��fŮ�Q��36-��/��א����2U�����q~K�ۄ
����y��&�?�(u�6�(?���b��|�E�/�p��m7���y����1�A��N@�A�?E�h�����Wd�s0%������ю�T ��*,��Yhi���gJ�4��y_Y�ޯ�,��������7��>��G�t�>��a��F�����c?�L��Ɩ��舯u�۾��6� V6�gh~>A�!3�
73�h�Ʊ��"�v��8�f[�����1���k;<O7����`�_� ?B�Zi�8��ڊV	�3�]y��D�W¼���9J�Q�*����2�4ق$^��¸�a&}<�U�dŽ�;9x<o鐓j�ҳ�EB��=2��Z!���~��E�Y�B���=r�m�� �Ԉ��-�������V6I���W���3>������ S���x.Ղ?�U�I�o�H���h�ٙs�z��J�x;2�.�$
��\�*��DL��!/��#�Y	N?{v�l�hZ>{9{n9���*
�9K�W/�����t45�O�B\���	���6��D5��X�N���Epⅲ(Ŀ{oi�-��$�@�a�ȣ��_?Z�J��,�U�D$ޙX_������K�fe�jD?���X����KF�xu$R&�a�Z��D�����u�ex9R�� �X{�UE��ʫ����5��y�C� #�U@�{:�T�c���XQ���;�NTP'������V���+���aS"�i}Ie�6���q�3�gV�_>U��g7�����pk�(�K�,1�(N�8��X?-_{u^T��e�s�?���s�t�~�W�`W{X$��B�X� p��j��I2�����nAx fC�8o��R/�gW�F`u����?YN ����k�� ݞ�B�[E�)�ʆ	/ρv>�L�n� ���耠O��8/��!��ה�����tR��JE�f��5�h�b��<�fѥ�"���Fb/,d&�P�~T�0'}�D��	��v`�z�hm�?ehD�Qӎ0�Oe׻	+�8K����K��[�v�-׹@�hՕ�����Ro3_{[ı�?���n�[�!�p�^��=f�N\_�Tc���0�{�RB�&�FxS�W�8���h{��W��6��G�B0��ׁ�l���>/�R�c�$3��Q�Bj�omm�.ƥ�ҀY����5�Yݙ��!��e�mB���Ć��1�+/~�>�=����ϑ�*�2짃��Կ�����6J��z������`�e�,!�\��LZ�'��r4�������_�x�����KW�D�"vz���i!�2��/ae���JaX������EIA�Y��̍79���o'�qo��O��!���n��K��s^�SL-*�"�3��,��	������JDg�V��E��3>���0]���$���v�}�!T�av�ǕLu�֕��-L�V�1�����I�%�\M�Z�?��Q	�\'����Y���^���D���oV�y�`~�����i��NȭzG�!�~�5'OG ���Ak5�ԥe�~�2.<iL�9���\�RBJ�C���k���NtM]�Z%5�'c���F!y�xzC���2'u�C�����,�d�R�QSs���;#��sjq�N�_Q�T&�vUO�=� �c��5E碿��Ǆ���b���������+Ĺer�)I�����J�s��i���lX7��xӎ����0Kl�/	�(�>
�"�_D9������$�/�E��ux(S�UQeGT�B�:��-�HiKU�N�:�(��)x��<�D�c�T����2�����u�}9�����Y��g�o���C�����g�t5}�MS�J�;�e���֥��0Rک���^$�8�.	��JY[�>����~W,.G��X��9�OU�l��5TQ����i#A�'�HD^��|IK���i1�ZD�V�?ֶ� X}��<sH���"M�B��w*��2"�nP:��yT�Z7}�i鴛�D�	 �oϢT��xPpb�-�N�	�$��H"Z�ѧ6��Y5��K���a����:0�~F�,�=0S0B��j�8��z�J��*������A�$�|�9L2��V�0޺�_mN��(���[���au�E����p����1F��u��x�4�����uŨ�w��!�a/LV�m!����q=�Ua��?Y�E���CiwN8�6=�z���Px͍!�Q�[ �y�o՟�t�4�A͝fuC�i��~yXU�S�:��w�Cw�pQt��B֎���)q�lY:�����[+�>hcG��/��^��~V�9�f}Ez�!�X䨌_��#W������ �>ʠ��μ䩇K����bc(�X��
H��������z}���0���1i9kQQ���葠�!0@E �p�G*��3���0�x�%b:Z���vtƅc7	nq��W��X�/�|�DP�.��#� $N�)�PN�Ř����X ��{g��}�>
RH]�Tk��)�h�~[��0�y}Fr�����s���Lܙ��A�fB'�d�D�5cF�\��O���ș��2¤*��I�yF}��u��e�N�H��ٰ�p+��"�;�θ�"�����*z\�,Bъ\�uN;-�6m,�K�<�Qiv�Ë��x.���r۞�"2����9�E��xwٺ�����7�=�4��u�(��$W���pzc��IPW�3�������ܛ�Z���^<�@���S��V��:��F޹�An�X���<i f�;Nu��"n�A[υ\	-���2��ȺEq�|�n'�k�*ɶ+U�?Q@��ɯ��������/'�@��`E�h��5W��G���--4�y���uUz����ZO(�&�J>��X}��Q�G��h7
]�K,��q���܆�v���g����h&#:ا��\b��W�ߣ��]?�]�񢉭�[�܎֞v�wī���U	�#U�O�kxm�W���6�,�px��'v���yl7�t��'�=峁��S�5(��5���v5`��^���y��)����W(ɛ���2��h_�-"E�vaz����YG�L��l{ڱ��Nm.���z�
SchIh,����䱟!�i��P�?���,��}�`��U&�ٿ��x����ȩ"��,��%��&|�z��Ƿ�b-���^^A�JD�	����DYul��#Ü..mR���F ��?FD�S�����e� ������ �i�ݞ��!_��"3�ӭ���9A�o�m5�~5�F0}�XA0���s2P<ѹ����3��ET��{\)q�w�-�1,��?8S����ɭ� pΚA7L\s,����� @E
�����~�����[Í9�v��i#�_�őY���Eb�M��y�;��ۯ��K���P]�9^˧�	%�]Vw��%����ߵ2nF?�����dS�5DE�U�����&�+p�*5��Gl����d{�[̘������mڭ�D�N�:�#�|SG��.#��{`��I�18X`��Ц�3� �Ȧ)�Y+tR��åI<ɦ��Q����o-e���)0d��]���T�^| ��tum֊ܭj7Щ�Bdu�7�ƚ�w�x�-,Ӻ�Bÿ�U�QtBOA�^�6�aN�l��Onx���`#@��ati�a�Rf��RLb�%��R����@4Ig4��i(J�z����9ګ�F��%c�ĲO&C�'^�,Q-$d�������G�����z���
q*X��������Fnˀ�}i��	��d��mi���4�<MvX��b�f��"�dy�B~ǲv�'9ľ�Rd�U3n��$&���;-_�;�/"K��FX�݆f��_��D#����=�p��Җ�2�^	��P�F��K>��R[�@0��F' z��ڪ�HP������݇��|�9�׈�h��8��,n��{,9��T�l$u���i!�k͒�o��wO+P���q��CdG{�PG(�P��������'�c�ʅ6��R<ᮇ2����kE]!�GD-�7�T�O!6���t���ى�h�X�$ֱ��ʗX��Y�xY����r���v��wRNԺ�Ѵ,��XOFۿ"���+/����u\�Dk���߸-����R�՚O���9����� �Y����*n��6�/:j�L�,���'��/޼���{��z�-q�ϱ�Q�Do�&���yk^���oҡ���z<�WQKi���R�"�W~�d@,��hx!�R���vϛp-���)vW���`:���?.��y�h
]�C��<�x�iI���FOG�����8.��wss�=WڬIe&��Y��aq��]h� 'p���d��4����1����_��ci�HhRNc�h�D��c^��l0s�[Bv]��t��`���W��Ս�ց$S�ƞv����2����]+����b�S]�Q9��O�d��lѬ��t�,R��))a���3pP�;W*'�Ù��K�-liH�P
�r�'H�����8�c�r.[� 
:Q �+_�51��,�����aE�O�Ď��ۡ��;G��vX�eb!�^F��	;���o`P>tI�M��ޞ�D�;��;8{&�v�b��<?���h�Q	j�6�b� �|RY�_̆8)�����v�v��	��^��C;�����U��$����7��|��� =�����~:2�VY�]ʧ�97���9_IlG�"�5������b�������P��k�e;�7��`�b^8���j��ۭ?s��烒���os��]`���]�j�̪�p?{w��-|���15�̆�XIO2�n��+��&Q�O�l[�����-�1�APD3��e�V=d�.d[��P���V�y�z����E�X�L'9��L�k I���;F��h�
d�(�t;�+��s$���$T��O��n�:RV���e����6�����[t�鮨�����[�h,AE����n���3��o>�j�3E_C/����$(��ys�Nv����}�O,O����ng?N~R=34q�HH�V޲�Y�RE�3��PR³x�q�M��B|�"���*?M�sl�?zQ���(�;���ql�FE���"n�J�.�6yG�mh	Rݘ��/_�=����G���99��A6��Ͽ��ǂ��y+p;��%����"�$T�м�҈���#��#��~8�_�3��./
����������F���O���'b.�ًwc�c:������Z�CE]�!�m���zÍ<^�DU�85��*���Z��r�3V¡+1GL���ք]��D2ԦUdtlYZ�IHZI**���1ۡ
~���>]R{	��xy��:�nqo1t�p]�A���sXl3�jE��q@P_�� dZ�l@�+�鶞� 0��]���'v�z���*{��BW������jE���|�����s�V��ۊU1(E�d:�s)�.��Χ̿��O5uu�,�Y|j�5�4}1%3 ��[k�{���zF���=����	�GOo	ѕ�x���P2�,�e�!�P�|���5�av��'e�=I��T�,m��~�'k��>����{��\i���EHa	�M��W��0��H�΂c4��3R$�u;.P�7��e��6g���@�8İ�AA?��'u� �/hc��E(�4��E>��Sh&���,6�:�}ź�}����oj���EU%������P����.F��`�Mt�M���˼�!����e�V��밧����Z���Ǚj��w�?{@B�ںk�8�=��Ug�Wg�qyU�t�Ѵ
�e>�_��٘^���b����7�wb��օ�ѷ�&����m����%�d�I)�m��u�f�4�$$5q����k��
�/���K�Ѱ���"u�^�ulB�>�@2�J����wc�/`�O=TO��tw���#j߹��	��ӌ���$�pqv��`�4}�۳��m<�;g=�M�`]Wyއ#��O���+|�PQ�AO��a����J:�(�J�ѓNK��`,PҎ&���"�\����Vf��k�[�<=�Tt6 ��m,�Z�d�i%0�w_W������]È�s���Lrb�50(�;����<[5i�%r�|��p��=t�O�{�K3�wH���:�'��9�L�r��+��Mc<�aC~˃���H�%�$Yc<n�����׍���n�HjL0��w��[?H���
s���|n���F��:��=T.ҥW��5H����_fm��2�?)^�?ڰ-����r#7R�.�3zq^J�{�w��0����4�,� vΌ�
��A�-��O�e��D]�׀��*����r����w�H�l��.�����O�^X�ځ�n#wV^~��v!��2x6~���0�&VE[���{�f�� U��\s�Xw�k�������y����l]���Tu@o�

pI�AY���$�%�XZ��/�XxJ&�D5�5�޶����[��B�X:Cx���yNE���`\����{� Bn�	���"���(!�e��x D.�R��8
/dh#0�-��2ʃ`��9�']�XG��U�j������4ЬB�����&P�\��ן��C�E��B�����G���_�~3��'��\�\���"�Ͳx���>�P.���.
j�����nA?�*:��y��Fd�lqtȪ/�rʅC�.h�w�������X�O��p�>Qw��)HE��4"�<<X�a�	��U�$���&��;�g�_r�����D�]�7D�Q���%�D:����1�=�G*�^x��EGs8�'ݙϕ��}�$��4����ˍ��^��ƸY"�bz���E�d�~� ��Z���b�[U�nr�E"?��Aȓ��:Y�� �cIxu���}����[u�����"�#0��F�@�:Ej��R���Ổ#�#��ڕK���=gJG2PpI��n��֟�<e�A�������,�����?RCER�2��U�$*P.ԺD��L�0�O������@J�_��9�����������������.%���ٞ-�M��� ���w,�y���Ehi���j�5����y�k��gk@ɍX���ŭ��`�F+�ڠ���,7nX��;U�~A>��tsS	$A��	Cj�" Zy�H����ZKL\����J�w����І�#FI���\7*6�o�cv]v�u��{����`���(�)j{��
{�l�@��F��
@$����]�F�$�Fή�
�����y�'9L������x#	��np��<��ܻ3˯^�l�Z(N:�5�D�\�#�I_s��
��k����D~�E*YfL2�3�7�iRiM7�R�Cs���l��}~F�GR�[�R�:���L�^45�=��h t����i�������2��&}����K?������JZ������.H���@G������:��/�iK0Μ��ba�q��o)�MJ]���{��A�m�͋��WF%jA��9o��2�6�ҳbܟ�Tf2 ���
�_��r�}W2�4��5��]w���՘��Q�zmB�����/�:��6b�2��U&TȍH��~c0�]����g���n���j�Y�)౮(/�KM`��W�����I�0�H�i/����k�'c�}�R�ӂB����o��P<�A%��
�b]��]h�ٱ��Ȭ�!���ґ[����ܛ��_��5�=
�D�)q���Z�vִ+������0�]K�;���@��,��Ya�r�^EB�|��##�*�.�|,}��>��(�E�,��SL�&V5,�B�)�W�#TO�O}��a�3>=?GL;�7�c�4���h0]ϯ��z��������Y���ѲZ������� �u-YSW����<�����YZAP�m�<�2z�Q��:6?'E�������ua�ﬖ�y���ึ�!u�畬�*M��S�c)��7U:��e�a	���,�#��<�`�|���u���a#�v�����	��du�g��֑VAx�}��X��_�w�bl{�.�U�B�3�isj$�I����tBf�7��դ�A�PX�g�Ck#l�^��[ ���!i�N9"�����^HȢDo�ܭ`����R�F����C�t>�ָ���C�\fRW���'��gklxC=��7�_�R���������+Ϋ(;�y�fH�!"C�aO ��@/z���I�O�C+F8���۪�tΜlU�/n׾��o:S�,�m�d���mU&_i= ����2��@tcsz�_��Cy�������.f�ة��=>�� �+�ΫA��>�ƁKQʦ�UZW�����%?�[��	������VVz9z=�>�a32��������n�*��:>T�f]b���J*�
Eٵ��7�*��,g@��;�r��$A�A2A*5�͖E�~׌CD�p�>�:��Y��k@fv0Q����,�[�Ӫ�Rl�72�S�J��z���Z?T/�.C���n�]�D�����j��0z��X
�C�"D�$ʴ��$C��/�&�G�2�*�a���_������a�����H�l9���_���F_�;5��o",8cL%�C�a���WK��b��>�l�����*�a��iH/���Um��aI�o�~b���� �����/�v�7էg1��,;E5�U�gif�.:�kC�Md^?7�(/tT��.���[�b7CN����H�3d~1�f!R�%��H��-7��a:D���+aF���.�u���C�XX2��m���������}rֽ�`�W�������ͫű����;�����{��V
��i�c�[+�M����*��3 9�B��W)m�+��k�)1\�o�`+�P�#mޜnp�mo
 KD��Wu�1�����P4�I�ӼL��b�+r�`ݸ1)���IyƑi�Gi��$V�nr5M������/#�â���nqW�g�����[*�����1o4�%:��-U���*4/�rӒ#wV�w���,�ri:��F����%Ǒ,��5R~��3)�����e�U9�̬X��K�xL���oM�+!�G���%�-f�d�ڡ4� (�"����=��O�ek��n�*�#���7&;�ۨ�E�D�p
=��17��K���ۦ +�:��|d�ƏR��X=��aK�hV�J��leٲ�Wq�ue�W�Mf�~���?|MA�O�
�|���o_�s��f���#��紮���p��1��4_&�x~LP��b�I>��s�b�S��Rۍ���Hօ�S>#|,3���vN� ��់���zE	5�� �5ԡ�f7��8���jY��T��@�wZd���!��t�$�R���>@ 2��\�W(����=y^��\��fw�)T4����H���}8�M@tX���\ثs`E�����n���s_�6i11S ���@�u!�%˕�U��Bf I�����=�P<��KQ̭>���H�3
�\��("�|�=�7ƙ�6d��\���~{�);��K�(G�t�G�m*��A$\r��}�YS+��z\�z,�2��x��3�b���܅d�����fmu��[\�?i��KwS.ޤ4�E�.{#ޯ��55�s�����t��aD�/I�۠ǟ��},�;P{�9X{�� �ϣ���!����i����6Pv}Q�GR��v��ڽ��{����x ]��ĥkN�M�@���\��x��x4_����nTZ,~��
��E�h�<�$cԫJ�i#��y�b�Z��_��V��eĎ��3X٥_���I�s�ćJ�0���*n�]hZG�u��0���s�<3�ʤ���J�B�&G�rG��ߩ_衴�s�6f�ٽ�f��φ�������x�c����AC[9^
�e��q8A�L�jk��MQbl\Ņ�L��D��S�'������;���p����YȄ4V�ٱTHi���:�>��p�^�������NQ �YH�R���j ��H|�R�����<6J�V�����G��R�APW�����Ea"�;p���ˇ!��P��҃Z��q=���U�N��p��c��j|����Cwߛ�2�L��&�06�)������| ㅭ�-�s�D h{y��%�z���YYȸH����A�hdx�,KS"����i����y�$B�mpd\����t�7�F��3z���p����ʠ1���I�鯷�x�8{O��d�H}Pv���� �1�r�p��8�W��������S�z�1)z,�˰Y�#}Y������JX�ҏ��L��"��E�4iX��I�K��S��Ss5o��t�a�c#7�kqh��t���ԪY#7A{���D�gP����o�d�9GXe;�9
��rnK{���n}M��JN��o��;TN��-2��E�o G��BF�T�x�CN��^��HE,���?ramA'���x�b&�D|�~~�m���g�.�I��y҅����py��� wK��%���
}�:�
s��=j���I\�gA����	G��:ߏ�2��n*�䌑{Q���-xޓg�N�����d�Ino�k��$�-����^4_ x{PQ҆��%�fD�#8%�>���(�u/?eV#�Jm�v6�d���#� É0����+�hm-���`�<�O$a �3B-25d������&�"\��O�R�x&���e�S=�6P}ʆ���ܜ	]���j��we�=aoe"�H�7<�g{D�n�<���k�����{JO�q#Ȟi9���8��ٰnw�)�Z���j�D�ͽ*���o�V�z�|��B��&�y%�׵��	���%F�a[�(�,}�X'g@�n�9�f�HD��;m�4�pC�WtOn.|�}��̲ηV�i�hP�EÝf�]��@�~B#�1OI_>�/jL �X�IO2�$4���~��^����}��o���>b�u��PS0�R����G��kOXg��|y\8��@�Lb�i�OsSΨ7�jf%�]F�Y9e�{���#൰1�����Mm�\+�B�c~�<+�3���q�Ӛ[Z��j��;7h1�Wk��$T��b����q�k���\x.\4q�a�RbN�R��"��� m�9����hvW�F����q,��:wr���W�ho��w�£�n�H�8ӆ0vM$�N]H�T$��q~���,B�a$7y���; qC$f�!<�k�.��$�a�1��Ï����r1�Ԑ mh|r�+i�>1/E�oչ�{�%z��(��n&�H�r�8X
N
W�m�6���P���7�QN�:*w�[[5)���u�xg������^�\o��_iC�٣��*^������a��t�N��J�D$�Z��~�"52�THe�/wM%��z"s,_4�����E���c������=-�N�|{�L��5�:h����؎Ϝ���nO\Q��Q�,�qe���)P�hfHVm�jRƱ=*[�m
	���&��%���+��'ȵɣ�ԉ�;��QN�a��	����5W����徠5@���/�8�Y� ��o���<�*}�H�k�����;bR�oˏ[����̌�\H���Bt�{�s��Q4�� /ԏ�-���w�ߤ�Y�X�ԥ� 퇫&jY���kn��4_N�tw�J[*�DL�
���oZ��������������xCs�s����i'w_�q���~�%���j��H��qy�K����Z�n>�_K����g8�]5�]i��\e\�u����K^�4	E"r�F�c�_��Pe4�����h�lY�t���@f�)� w�6��ZYBhŴƀ��8蕃��z�gfU����.
ЭT������o�H��h�.������]����x�W�O	��t����E�!��=��X��!AE�y%��]�>����ð�@�� 8�*_�*��+�%�:�"�x���&�u6�O#i���/t`�X�a�/s$���� e4�LT�	5l�Y٥D׮��#��z
��8�#�t1�m�P���IBE�.�\@vPn�a�p%���FU�7\���=�e��3����j�a1��ZU:���O����p�EZC�O�xܓ&�O��i7Z��5D&�ax���m�-K_Ar׮����M�E�	1P,��H�Ȝ�D vh��<hdfO�F���}ջ�G���*<��5��D��7�TI״���4�����.�.�x&��.6�]i*�� F���/
U�q���^"�@%��1��j:���0���i�����\-���Mn��N�I��\�"��L��髹%K����Eّ�p�P�O���
	,�#�v���m����S6Ճ��$�F�<E}o����5?��^~��UB�1�B��l�P_����	3#�,��˅�����7�����)�Y �m��YE�!*S��ᒘU���
{.�^k���t){�����d"�=&e� �O��b~M��5���^���$ȃ_���tqɉ{�O�PW����q�׼7d��90M���#���!�P��?�}d�����<�]3ëR�9�&| x� �
�|���c�8@�i6Fa�(Ş���Ћ�4wǋ�X�G�3s���ve�\_w��;?��w�~��@Ӊ���m��5����b+I������x�y��
�L9ɀ�a|ɕ^oO~΀/~j;��aeЖ��p���~��a���(�{���c�u�O+L��hؼ\bO]-@�1���+à���%(52��ia8׈qQ��`��G�׏\�!1��3� \Aw�Ǘm����}�cL�a>�U�+u:ʩ,�;u9��6�k��S�yCO��3W�ǈ�)vCA5�"�H�����ۦ 7c"M�h���+���Rb��%V5.��2t\I��,9�
:�ˇ8���ХG
�d`��_�y�dK��)��E^s�ΎU��`9V��B�!�<	=,�fTG�=�h^���X�&OIR�Ā��{� i��5���9}��՝��7*�Kt��+<�Ws��پڐd>�]��д��i���iU����_��͇�u
�m����U$,��{K��Z��A�#�ِi�d����(8�GY,�4;O՜�M ��s�Wur�����XMa���+t�_I��5���tI�	���������{UI�8vt�¬�g�fIT\����x^���!�y���v;�x{�
ϟ�69v%�e_�||5� M���gP��&�g�ܖu �x$����n�^�)��J����
��aD��nJy�F��x�og�W�N9����ɥ���^����~���aBؕ�}ߨ�>AM��6�o��2�-�_p���C�&`Kt�<!z�!��!\�X�]���q��[:�m95��e4��ʡ5��g��M엜]���Md�և��;è���5��X�ҟƣ{�sbW�t�m�:�b�άa�*H&����8qH����,�4�8�f������[u�\|!iN~��)��?�;9�-,��\ǹI{xd�rƉ
�	~�������1�&�Y)�vܘ&3�Htu�h���"#�@*n"�=��B���\6�f:$ZRn��w��Tf�5�mA'�^$��>�(n���Z$��x��Vb��x#��7�����x
�y�JX��im���-Յ��$�|�����GF�γ��XM���,ߑk!\���ڇ��aޯ�`�ڻѢ4�e
v��n¿E�5Y��jzG���:|�＠�-�a�*��[�������d*�t��G棙�)2����2��谒[���W����Q�O>�\��8<d;�+%���Q���~�x��e�Bz��'���ݧ~uI	�(�8��"A*�z����`��Mh�
�����DU�]�n(�F�2��z�UG\����+�?>�"Tk5X�(hw�m����[��a��:`��+���e���slNFA�&崔o�fq���@�\A�������'.7)�B�����J�>±���>vuRHP`c�WXH9pC�Mڣ�^�[��I�o���)왘пhVSy�12�uF%:{�������4T]^�W.$��IL����ID�/�Գɼͽ�ʪ���&<���#�YJN������o��;�#�����/��Y�����g~�����V�/���X/B�v�����E����i������(I	=)��<���W�'��h�����$�.n��2�2f����TSZ��
֣����c��?}D���d�����y��������A^�x�eD�D����g�����SG��E׊�w�$Nl
P��/��w�%]_�T������$���Xp��;Ǳ���N�Vб��)O���҇]fIޭe	�i����lғ��0?�ap�a�gݍ��f_h��/<���z�i�J�{
���ÿz#�ha���u]�D�'�Ef��L��3��\
 ͺ�3�Ǻ�	�{EO�}e�%��x�����N�k6A�0������%f�'{RtRm�b-ՠ��U2�
��

0!�%t����LC�D]�1Ð�z����-;eFG!�4{�3Z����-�z��N����I�����{��K���!J��|�O�n�ܴ���k�C��H����x��6���D&�i��^G.�s.�p�͗ǘ(�Í*�"�7w\���pW���w��@pca�Y���ᛰ����8R�P¯�!\��˔7���9$��=m�ˊ�J��~�b-�LwÏ��"��~�(�5K��mI<�L��%����"]Tr�d��k(W�&k��QԦZn����q������=��J0���{0<Q��;��]H����uZ	U�X�OL����GG��y.�D_UT0���c��Z��"^��W��L�M���L���w��*W+�Hx�s������ �/{�=fr x���>U���5:qIxU���c�!*."	�8'|�^�^=�s�?@�c��0�s$G�{�XvK�����[�3��+�.����Fz�.^Sh��V�!��zD���bYĲ×6���<"���~L'��+#�[B��R��W.+������Tx>�X�'�����|PY쉣|Y{Ѻ�Ma����`ʽ�"9_��&�0���>��оip��@�r���޴�b��	��m7�t�����R`ŧ�lVŜԎ��e�+��o���+��nVJӊ'��M����b��MU�yl.�5�>C�H��E��84Έ�h7�[�Z���i[�9���M?$�4���M�ǋ��$1>s�������#�A���}4�j��C0���"ԁ/:����Z��@���%L�z��h��5�l�����Lz���u���"��\�\��hUu���\~ȭ^���φ��0u�ã�~��P������M 7����6G��M���@]�������س��*n�!��,fىɨ�_�O9�Ctaxo�����P7�,'ֶ�:�8�@�x0ai�T}6���9�KY��?ʹ"W��k��u�1��8��;���nS�+��E�-�Ӈ��v�\8jw>�4�L�?`���?~�$���7���|8�\�?�v�z�L��
XX�QG��-���DN�K�\;��6�p�/�$�E��nV��	j8f��j�	�Pq����dL���'�|&sD��N��������I	_��C��4�z4ʃ7OȍD)�d�\��ۑ��Q/[��
dR�e\�7+ܵWu"��Z�U�|�I_���z$�'�'��Jo"�}�'�xrw��Km���F���s��;�Đ|(�c#�z�������@~�r��AR��8��⻏�Y�8�8e��'M�{L�)w����Y������M��X�ä^]��ے'�ŤQ)w�M�\��fۜ���^fw�?Mʏ:��h&^�bf�:j�`}�t���*_���-�:G����;���1�M~��T�jܥV5G�5�rLfP�,_�"l�a�;j݅��M�8>ı�D�r����jv>�Y^z�S��B3ΘF��DM80�K��Ē�[R,�q��#([�y~�%1����g���#7Ô�,�����Kd��y"��D��J�~�f�)���+��k�X< m<0E�/?7�%�Ҫp
}!����+�����	�,��2%S�t�ms�h��<
`)>����1W��/��1���ע/x#���`�u��m�ş�t�0��$t�R�3��+d�~t7_��#��m(�����_����8��d9�~z�"��ɹ��!g��.�bkL7��꠲�|��2��������}���>W/D5�����<T�R,Y�I��&J��gъav�� >��2��>��n?[��Q��6|�`�Y�O�+�WW����R��#�ݪ�L�@����m��n�P��
�#n�x�ͤչ.��4s��skJŋ�����N~:<�բ0���6
:Q6��=��Qq��B���]þ��a��֦vX/�����G��H������	��\�A쟲4s�$3��Toc-�iМH<k/	��/��r�I����k�h%��/:�v���0]�¤�.�(�nɄ�hv��g���p���M������B1ؔ�@��;�>�#��μ����Md� �+̐v�<hiЈ2�ݤ
K��|3�<��Ip���\z���aQs�]VS�<=��k�'a�tB94��|�Imp/���-�3!�EN����Kɚ���|a�!��W�!W<P�� �bw�L��uM���ᕪ/i�����aZr܏z�:�p ?[�u�]gJ6�E�	�{CC����r6�Ę���>��Q�Ch@h*֬2@����y;��S���l���\�q<<rv�)��r��,|���������0O������Z~�J���U��m-���l����R��冯�ہz$�[;T�r�����\���b�2e��z��fo#��MY/gu�"AX��h���s���@c�yD���L��DU��P�~��x�74�L�����^y��o��4@*��u[Z��4�;'|� ���!v�]��d�י�G�R�W��� �����~��+ñ����ͣ�As�kijr�W�.��KT���Tz�<�vyQ1NYtRz�S���>���q{�����,�z�y#oR�y�N��Nh�Ǳ� o(5L��{!�dE�j�i.�|�sp�%�p�8+,Iӯv����"�5�$4>Yk&}5҈|3 9�,*��>�a�.�V6-���Q�M:��Ȟ:NhP(4��5Y�s��d�����b��?C\X$��m7(�_c$�J�G��L	��G
�Q*�X�zy��r�l�	��s<Q��r���f���땨K��T)�wŉ ��]�wk.�&�{^+�W��8������
߶9g|�X�xS�)�[0TūȀ��9B:�-�4��MmR��ҽ �8��"uRv42�խZ��8���yjU��I��u��Oca����>���ڶܮ�_��֑."_��b��\���S��W櫃xd���}��[��F�6�s��yA&S�0	uMLȣ�ҿ��?e	Y�ZWa3)B��c��5F`r鶖��iY?]��7Hw��B�(
;i5���tE�)�?p3����$�}��n�@������1����=����(B�O���yΕui��Bh�l)%�kQ;()�J�f��xǢ�:�͊�N��EӋ��F$ќ<�lƿ@�h��#����w*�2w���f�H�r��,��B�<	���s���7z.���{H�;�pQ8[<�h�`^������k�;�jn�v$�Q�,�2���>���#$X�羆�R@��D��`���	,`Q�Lk�+�	�6/�@n�覍�j�o�3�j�:�����Tw��ƭ1M:�m��6ه�UǴ�p��ߗ�Ŕ��(��O�/3����;Z��W���f��U��ĭ��ځj���.-��Lzvr�X0z�]lKD��F<��(��M��5Ԃ���Tۚ�4R�D1���q�����7���f��u/�
�#��z����#S�eJ4�=ڄ��5�)%��у�d���U���x�ps=��~צ��*���d��U���͒2�_�z�>S $U���/;��y�����G�a����ޠ0��y�����i�d������_%_8|s�"n���{�/��b�y��B.��}���$�M��!
Q�1J��e�nӎԏ���u͘��@��"�5�;sp$� `��2~����Gg�XC>%a%�@!3��P�''�s�@:Iљ'{q�?*s,���5�Q^<��F���
�1e����ً�D�݉��@�P�����n8���" A<I#�a����9tʹ-}�X)�0�U�ǷY� b[�՞	"U@鋬�q��I!�_�ӗ��g����H^�.TU�.:�C0�VB9�G
[fE�7ӱ��zIz3+`����+<p�%0h�瓾~���mq�`A�w�]
�Pˍ �{���:���E�l���8r���W�3|�(aa�ᚾ��ܣbd/�S�r�qDp
A�iҨ�G�_ ��U�Y4ps���.j��X�D����2�`>��bN��u�����WF� iW�ȕ7��lj�>�D�U�M�?e���������88d��.���-S���6E�qp�S����!\���)��W$L�'1��0�B>��A8؁��czl��y��*�>�� Gq5ni��Nִ���VP���9qX
?�z"A�h���������OX�p�/X���HӪ�?���h���1���=\����_�	S{���=�yrJ�c���wR5Z�Ju��-|?�����gQ��ЊB����lGY�5����g�8 ����<�@�]�3B���Q9�AT5��*KS�y��U�f5����A�a-!�@;{�5o�7����?c�hEAk|^��]�=�E�V��H�R��R.��hE_;^�o)�*��(%P��-R��?�u	�K٥�S�g0i��/c��l�3��x� �
Ƿ|
��c�����-�ύM.x�թ-@�3$�gùtth�ZӮ�����=ҩ����Dͬ�Z	���і��(<��;��ib�]|�ɇ��� OD�Y���.�nQQ�J('��g(j=�����u*e�7��p�5�)��j���}&�C��΢���d�&���nS��a�6�- �6��Z�RH������˖�4\ǟ�jG\ +�I�L!JO1��?⍄$W�L�28ٿ����rwnr+���0}X-���I��1��ћB̵K
\���_�}h(�c�����0E��$^����r�b0s$��p�D��xҌ�n�o�6�q�"5聃�?�ubKa�O[�J���Y"|_Ipw; ���UXt����.� HT�f|���VЛ�ϧ�ͫT�8���ֶ�RE�I�G���i���:@ty{;ĥ�i����׽rO)21R�8�/�u��0����("�V[B,'"���`�ҝN3g�"�"��s�y�|S��u���!���eiT�l��4$����7�@
3��N0�O��&�"�'�!�/9�����B\�ML.�	��A��e���0����p�#ȽVT�A��=��>��&h|�dpl�k�7Ҧ�STP��Q�&uz����dt��e�Ÿ�HH�\�,�kaPC�O��hmHcSZ$����F�q����m�K�HpW{�4��pd:����y�+��q��6�c2u�c�J@߰/��o���4��ߙ@�~(	�}'q����D������luaOh�@��f(==���D7#7�[]�:��� ���lRx��"�^eu�� �B�op%���rDzDj��)�����k$�?܍�N��:.��VXx����҈������g�q���Xrs�}
Ъ�:p���6��>+X����B ozD�y�3����<r�kh��g"�c���.R�/;�$�X]b�J��c����"�����B�%�tL��H�i]?+N6��g�[;�E�6���+5i��[[�|'w�|nFͅw���u͉�șs��]�´�8߭Jy�v[�<�E��zw�lK��3��Զ���4���5���:�,jɨu�=v��,��,�h�o
�����,�������~=1u��P��߸y�8$2���~��fȢ�@����t{��2��S��oɱv������������%-�ڙM;)��M��9�m�.|i�^�t�aVl��挋:���U��\��7��}ٖ����6�s��G��O��,#���a<�����@�󇚵��J/x��RE4	R�)��P΀���A
-n�IT=��ݎ�./�Ay5�(�Y)�i��S�1�^[o>�@ڂ�˵�z,�OpWa�L96�|�կJ��a�c�m��>)�z�j���!�f뾳8!�K�H�����k@\5��>,��ih*'�����b]F���A
\N1.�����N�0҂*����.�5�(k�W4,�oh,½�Q�^��f�놝�h�4�:I鷢�y�ɦm���	�@ �b���E%6��g�!L�=�Ù'Ǘr�B_�!�z11�@k ZV���;*$X�UHFe��[�sD������1Hm�k�Zm�#�ħ�r���5[f�*]�'�>������� A=��i��sSsѪ��mM땑����f2�U�T1ƠZ����6N����SD�t�"�����b�WM�y�9�e��7F�����G1z��z�NZ�.��]RFf%:��m&޶���~�"^-����Z�׌��6�{�����c��2dO߯�b�<x�hK�)O��i�]���9��_�I<>��P�^m��JC�:�3�}�<�6���\���S#YkY���wf ���FV�ZHU�]`�)���^K��\���pג��g��_�)>\g���tz��l���6�6�^ER��/�g���C����h�ݘ�h&F�̪��Tv��R�w����b�plo0j7L��4�"��d��F�������W@����Tô�ل�0U)�� �3aU�R/���#)��I�Bu��`�����$Oȯ�^p�d�k�3�Ҕ�@�9j6�D�0����d8�_�C+\�����x^�],�(���{�)a����MF������w�S�λ���-	�U⚩z�8� �Ii�/=dE�^e{XG�YI�I����R��y�!��jh��W}jP�\/�P��]���!%4�5��˓���8Ȇ̽>ڵ���YS��Q�n8Yhl#R�^��B�d���9����[���G��~�`�p����#Y���˵r�ٓ�Q���F���5���E�3��^_$"��+��m�OЎ�$�e&�1�Y� �ˁ)ّ˫�cà�p����u�S�Y1���]adք�)!����;=L�^�l����S�����H�!da��p��kا��8F�ۯǨ���Y0�}ի��z�-N�Nc���K���F��(������>���kE4������}�"����s�P�r='����c^�f�`m�DQn�񛢋p�����0�$�<�d�0�~���7���'uP�������yXcM
��z�_ ��J�r�0�߈���A�rc"I'<~�{؍IN��h(w�b���!n��I$�kn5?C����x�p�#Ȧʈ )�`��gϰG'.�=L�1����|H@��<Mx�w�<���l�^@�.���	b;fPZ'�i�^Y8�QJ��Y�����L�p���1}r�� }[rѩ}}"*�&�R�@�Ž�F�ZF�'=�R�6�o$o� J�
�J{��5!NhV�xࣗ7�?��Yﱫ�t ��C9��L.c����)�nկ��}����ls���Y��7�i�ю���t:|KjB�|k�5g�����U׸��w���	:h���Z%GPч_�EIZ���'В0P ��}襄���}/�B�W,��4�+�\Od}�W��+#
��UT_-;I�)���v_Ϲ��x�	�4 C�.׸�(�����/rs8?��,*�N�����M+�v��-�4��m���tP��������^FySk�	�"�f(���S�.�^��J��ց�3egv�M�9��'hy!'<i�F�_���s����0~�G:�~��a{�Ȃn�W�=��<Ⱥڻ]��-�@���^�͂�F��M�����[Э�
��Q`��U�|�ܦw�ݿ�<��	>D�DhS�E���)�n�	
$�V�I�\ocz�o't���Sܴ���HMF6D�y.^A9��I�~P�#��~�pL:���Z[u�M;I�9�Ի��}A~����6#?Iϋ���V��\lL�\�D[��[�:K{���qqC��ʙ�ޫ�������uI�5����M��~�2D �����8�m�M�Ȑ���Aܿ{��.c�0`7�	� �X��ϔ?�"c��NG�6�)����dNs�|��Hp�`մ�f	��ޤGe�tj/=hR��.��=_5�1zP��+��ì�.��5O}�G�P8I�]z�sO�)< ��M*��瑗P�G+�n�Tی�~_.�K��vФLO@"g�]c�5v�Nݝ��,Xb�J��tOc��Z�k��q��O�_���0k)c���nE�ɰ�����峯|��a�q��������n
�ۂb����L`xȟC�uI���|2KI%�l���z|���C��]ʦ�u]2��W�f!��_f-:T���\��:_#Z�O����L��[����`[-��~���Pg�*=���K3��ŵ�OE;G�l�3* ɷ�Ě��Ҿ�-��
���4b��Q��*�x�1~m�W��#Em�x�6D؊���Ъ82_V�Ml\W}6NK�9%lo��]?�ܨf��[�M]yk��[4b)����Fѻ�]����+�h�L�8����6�1��[&��
:hJ�R�~�1e��a���Ǩ�7nN/eO3�p��J�|�vk�;��k�Ik���R��Yrr��j��viӯ��Ο6��1��KD��lߝ�Q��)������c7q��j;�÷�?��̉K���PT�1�m�'�[�I U�m�0w�4� mV�=K{�R�y~��i�wS����л^޺b=�^:��&�i1'3�քpv�s�p���e?�Vs!��'L,Yc(Y4pՐ�?�s	��\�����)@\X�!�^�g���%����=eSk��j�q��{jHu�%nQXP��'U@5	�-�1BC�^�#��_���¾A͆���Q4�;���!l@����T՗���Uڷ��U��~�!ߧ�(��8a�����h��[��;]�[d�]`h:A=�{�B�s�TT���hqj�L`o6\Cy��2&�����
3w��.>K;��?�̿��p>��\D�:�:�N�2�c��	������	7�<���@����B�
��Y�n=m̳�P����yV���3��q��W��ެ���)�L�G�6H���L�*�zZj��i6����_aV�5����[sѵ��u�n��8Դ ���1	zrrFn�������{_8��7�`dB�;��Ƕ�-d95>�_��E�7��ލX�Z���b3 s}�M-*���-�9r%�~�^㿉�V���u)~��z{'Fr�>�[B�q}��������0����澕�E�+�r��p4�2����킐6X0XZi�����a(3Z����&�WbmP�93��$��dx�%�P73 {�A� �l|��c��	y�%��Q���1��-#��9�`��K�����Z0��}��~�0�n�.�I*��%�F�-�f�Ih~��I9�4w�
<Yitv��>�id �9㼡���?5l��'�&;xD Ϛ�0x��䵥���!��
I|��6	Kl�#\�F��6���2\B�II���L�?V��Nθ��M_�3�|�D>b��^ �z��^H%m���Iq�@�..VBW�E�F 	�����g��B��F���^#�ImdhG�;S~nv���&��s|_��d��q �/�F��Dؠ������s'mm4ub,��A����<�$��l�޳�dLȋK�*���@r4qʈ�π���W�A�dq�!c�@�.�t��\��֮����-B���Urn�Ws����ګ�)�,�(>�	 ��f�����iIǝA�,�ۼ�t�huFM�4h���9mʢŲ���zk���cZ��q�鼦��\m{e �Y1���_ ����\q������~�Y���Q�,�@$o:*���d��޶i}2=�I��7��#�no�1��ff�ҜXC�8i��28����i���m{,�������}C �)z�}ˇ���mk�'���S�y�E�α�.c����m�Y�J��R�T�;�#YM���u��x���^� goJ k���Po� Sl8��@���(ji{4�"�n
`����{?�M`d��+;�g0k8RC�I�t��l[��ھP�T+��#0*��H�]�v�x�`Cu�T�H$4��9���V0/�~�� ��Wc���+��*��EK�h������A���)��3�R�(z����@Ƹ��޺0>�c�(�u 
c�k�@��z�39k계�B�_�E�88�Jv�=2���4B|ژ�d]9G��!��%\J��S�c&c�0�Ȟ$M�=�<��I����m��޳mo��$[#O�$їL�6#r  Ly�����`�uk�������S9$���@4��>����)�JБ�1:��+�hZ F�l�=��?V�����#�@��%�#D;�Q�ޝ#JO���	d�q�$`��>��+d��g��?Bj*:�7#d[B�5CW�rK��GK��B�tv��-�����>� .�9㵫Y�x�Ά�u�1���Ƒ~!{�mNs��|��	�0��<1���ͯ5M8���e���+_羣ݽ�݃�{@U�Zz̫я��#��7tǢT�J�!�Í\թu��1�>���<�N!�YV:{F�A?h}��C��V��F+�:�T88u1��I��zs�Xs���QIu�����Ar�U���J����D�Iҏ��?X���u��SʜrVDP7�PӁ1�4I@��J^�Xf=�DZ8��B��Z<��zLI��<�Ӯ�&�2���UZ-����ϴn�!�k8��0<��ameQ-��=�JIq.r�e���;j���}6�k8�XD�ZXD�$j�@{�C�kтMD���R�AaX�ld��T0'պ� 'k�5��hFV���|��n��\�i�֊�Pg�;���XB�9����L��6�&��!�a꜊�=�O�q4�͂�I`��G��VS�39�á~��f��J�d�\y��&?Ma�Nk����2�c1��
i�+q�/�^_�7�j��'�����>|@`�����F}$?)
+�D��`����-#�l6�5t1NB��[� :'��X��;�l6�ASq(k��6�C�2����������-��t�0����<�bSh�	��T-��3��<�_��H�5S���8\m�j�y%�
�}��?�/��|��`afYE���UΒkw�d���Ϳ���g��/>�qB�K�J��*�i�ߛb7���!�~��!pҡ?Y,\�W]p�#Y�ak����e!i�ԗ�:��uք"T�@��l�K���e�5/"��E��B��2�j�����H�O\���p(�y��W�Y�Ͷ�G�:@Mc�,�;��)g?v� �Vev��й:!��n�B�Om�Q nBrH�	b���@�WE߸g_1CI?�ЊR��E6���Ua��
�M�C�P�|̎��%���B����.�:�'~�(ȵ�m��u��j~U�"l���]�R]d�R��ͱf�Y_T��������TX%f�����Fy������s
W2:�.� }��~�=�dg������ʧ_js� �u�Ѹ�d���|𒣿��%6��0;�b�@z6ps�������|a���6���pA�RQYU��x�q�f��(AnZemJw��Z~��j?�[���GE �i�l��n2Z��I�,3���mB�-���[�L7LM���zd�ў;	}9K�Iǒz���m��/%�PNƝE��Ei:J�Y�?���^1TՑ�y �j���}��6�s�L�k�AY�/!5�XP�j�">0z8���7�.Y5 ^m��V�wB��3��#��:�U��T�ٝq��B�y�������ķVp��l]ĥ<Z}0����s^�+.�����v4E�D��W ��u%5��-9�u�(���<g�2�Ι1�?ȡ�q�E���Y��(܎�s0,�E`x�3<��ן�7� �*8'��su�@�ec3�T�_�m�f��1i�ڢ�a�!?T<�j�{��k��0;ԅ��;9f�@A�q�x	�0���\(*�����p��k�w�d��ݞE�������!z5w�!��$��χ����6�O˷Yt�^�1b���X�U]��`w�4�|*6�������;���2�u�P�Ҡ�F��_9Qq��b���b/] ��7g�
��{#� �1<��R+~����Bc�.
]ؒ���@�:/�QnU��8�"�F�̲3x��G+W�f��]U6�_P ��0����N'���3�\X�*X�F��lbķH�3�b�F�Ȉ��^{W�L�8�B�2��2o�����~t��&yz=�����џ�!%F��=��^�P>%,�d�Ċ�`oWq���n��.�U�G���ռ+�sU�`���Y�L�O@Ef�q����
�\*�5�誵�޵��c�̗�~ۿcFÏ��Ek�憨�d�M~�O#�w�[}w.���>�
yv�v�	=\d�ێ��ܗ �����+���&,	����S��B@:�5�5�¦�Զ�n!Հ�5�t= ؙި =�-��ߜj�"�
L�G�\�&D,�֧89*��oD���V�{�˵yAs��р�!^��a.*I��,���[���.D��a�U%uH��	�NPd��Sb�/+t��"Z���R��hP�����&أ|4�����@ֹ��䆽��a��<]��{|������P~V\'�	��C��m�k�'�J/���VL�˷s��
����[{���uHIwi����C��Z�{Z�E}��cL`���Eʕ�n�u�u��8¯K/�ܼo��n���QӰȚmCw2��@�
��UHz����0r#b�j��Ne��9� ����ǏbݍЦiH#��A�L�r�������+�0=�s���h�m��D�����V���Wu���tQ� E�ex�m���ש�o���Υ5`ru���.���74f!,]藙��v���S����uе������lg�w[�M��)�����u7���`�[f��w笉�@�Yo0�w�`2e�"�=3/$&�7���d��%�h��}����^v����L��R�Y�~��t��v�u��2
�RVL����\�h�e�C��f� �fաH�h����Jq	�x�p�]&*2��p�NH`�L�)Lڗ9F���`;\�����D�G��7k/�#$�p���D��}���w�H��� �G��P��s`�k�.��VN��~�4bR�����3���J��/����zS إӤ/�^�I'��߄�e�\�q�ti5nIь-"jس�7��=�35�R>��MO¦V�VyPM];ڃ�'�Cr�HD���~u�:�\�ؔB#��o���f��C�q�;@ފrɏ41c�R����#�2�2�n^?�f}�l�f�p��qQd<��p�i�hb՘����/Dg*���;�W6�I��f�+�R��@���X�})HRP\����kX/���q��� ���fBժ�;5z�=<���`ӓ��h�+�ka�F+�����Q�ӛ6�.�ֲ�rk���b�$(���龺�3�eZX<�b�U�i5������c��j¸_nF�������p|���u��Jc�8uMMv�c��*~>���iU��9��p��Ht�<t�Uj�� ��syU-Y����7��"�Y����2&v��Y�_Ct)��M�F�ܓy��Q���l�C[�"f������Ȉ�2��l�¦̸#g����� cX��r�
#��%�;ȼN~���D�7J4W����u�����$͹^a
���8}���+ʉ�DP ���g��u�M���*ci���ޯɳ�r�o��v�
����RH뒻�T۟�,ڔ��.Sq�7�lm!D$�E~�����k�R�+�\�P�]6x�{P�n�����?��I>���#��vyLt��%�#�܎���"K �)5���N��|OO�C�o�+B�K�Cg�G�>V�Q��)����ĜX,P�~0{e���/\t��
�R�s����NؔU�P�=��� xk@GktN������S�	J����יd[8qz^�t�>1Hņ5��S�E�6d�q��<�E�U6��W|;O�(���϶�(o6.0����H�#�,ᝇ�l�՝7�<�Y
k����Goe$H�x^����<��-�s�	"����<�/�\��pu�CORw�}��b2zr��t�ߣޛ��GaG����ϕo�j`��R��8&i�۵�0=g�m��ك��e���`���?���$m~Y�.�:��&6*(oL}EDb�7w����r��dt����t��q,l����#�O%Q&�\P��U�v�WShp�-!��mˢ�?H�KlI����\a��x�ͯ�t��T�<�k����~cZM�w}��-^�g�f�@���߶b0��; ����D�UocE%��A�	�2�σ�&h0��@�Oˑ�T�`�Po9{&;�l��o���J�Jn9�\*	���W���ˁ��
��
JAeO҂�AvR������0ST����5�-�5pH�u�S�$�� ���O�p��V�L�z��]���]�{[-c�"�$}}��ή��F �Y�$�TC/�v~�ʭ�tLƍCYgy��o�z(�|��5>����u���Z���B=�����!��+���.�(W�#"��?Q�v��A֗���/���;�݈fڭ�M�a�*-D�0�W��+$��։ �)�бe*�Lk�S�e���A]2��s� ;BU�����s��d��Wt��XPNQ<<���f�x>���制X@YO�܌hݛE�ra9}렜E��M/���ݥr�`��ۄa�yb42L�MS��A(}|��H�_�tO��g�n��H�X���!���4LR&�����]��^F-9�{L�	��ZE�k�QeS��FF{�|�v�2*$
2#j eWp��̫G��?����� ���PR˹;;?m�侅�\�N���]�əH@y�,�Hp�(�u�r�q�B�X2�3�0����Bz;��R�Mfa���ꅠ�]�i���MuZ��ZMt;�S�,�W:u��Bޱ���c��4c��=�[�,:(�+�DE�G��C�9X]N;�����~�j`:4��w�;�`��W
�Q�#�&N�=�(��,�C\1�m܊�� �C!N}/�'�} ��̞2'�+���~M���/�M&Rž���3?PމA����
�&��E*�Z��y����Oϰ�iR:�C��soy��b�04 ��e؇�SO�9�����m�q���
��:]W�y���^�p��cVr݉4���O�j(p�#AU��;c��j���xT���NJ�?G����q�b=����}y2�	M�B�R'ڥA;��e3�-�&(��Ub�zV�=�9��mρ��d5N�#q���ۭ����hh{���(�;�������7�p D�17���f��b���א�\g��̋�����T��`(#��S���<>}+���T콑w��if@��|�N`+7qHS�}R���^�<sj̗�KvE�����e�!Cj�����b�R����ҙ=��O����^���g�|("��vZ6�B�B���f[�=�����lǹ�����Ia4�bLv�^XE��l�.м;����3�#���dO|Q���:����6�UE��m%F�7r�
�%��>y�FO�W����/0�D_�_�Je0��P��$���R'���낣V9ѶL��Ϣ�b��*�&h1P3��Z�\8ƨܥ�6<{��^զ�]-j:�ᣪd&UmP�*\�O��dU�C�(�a�=7� m�G�#u�6�%dqM��h�׀/�|w�ה.%��:�Uӱ܉Z�0��)��Wh��e���Kz��S&i�bQ���8���F��>N�j��pZ���se�[��vD��V{�s!�}~��k���;��-6�h?�(��LF�����B����F5%8� �q�ǘ���Mu�W�=f�f�����9��1��F:}�D;�q���>�|M8޽'�dp�f?`��l�2�;���| TE
w|1�[(暫D����ዱ[���'�:�q3��>,���;�_PɃ�e:_�5]"�X���s^?�A=U�R�$�/�k�)�o�g�}��x��sH�e+7�K\�*1g٘��/�G��SEѽ����]Sy�P|��ª���S�����G�4А"�@MD':TJHy�:F�F�Q!+G7����Et��:\K���Y��X�a#
�g4xX�T:�۬��R� 
hu,�ev ��P1�	�k�����)
e�s9�4a���݋(�C�����*<E���Eb���C.z^1!�b3ػK���6���K�]gJ�'Vr\收�'�|�o&R��0�]�P�z�l��>��I7�ǵ�OHz���E��v&/�V�2�i�P����<�0j���~����,�Ƞ�Z4��S�%g�*�,
��s%�C�>/!<�e����G�K	��8t~u�z�;�>V��EP�����%Y�'R�����ܘ��@�L��HǞ��B!OZ�Z;Ҕ��+K��;�c�7���E0�u�$�4��6L�������G_\N�����GH#��l��SZªA8H���G5��H^$��t������k�גP�Å����H��������}�M��$
Fw������A�I�<��V%0��b5�}[Kp�~;g3�ZPa���9fk*Gi�I\���g���2�q�:V�}�ꐍ����D� �R`�y'6�����-�=�sK��ɖ�-_Q#|��r�ӓ�w�|��MN�ô��Z��wsfa�1k_�چ��l��;ػ����A�ڊ9,=If�B�</X�=A���J�Or����NPi���*����-������K�8�œ �9!��]I���kFP��&��D�7$U_�|!����8d��K��f+xT�L�X��v|�+��z$�l �U��En���D���s4@]��_��2�;S-�#�2�rG��ÊM�Z�UV��{_%܎�������J(~�I`$_�+�%	�R�p�?��4�1��M�%^h�I�ʹhW�~)�W^-H��e�ě��6r�M��B{X��M��O�p	�V�X��q��I��AP��Y�Y�x:%4#z�;b����q��e�tutƩ[j�҇�C��N��F[Y���Ѥ�͢��8�M��Kt�	?YК�ݔ&����=ܖ~���9[!�(�cN�f�mo7��q�~@9�(>�6�'L"7�v!��Dϩ�&�R�EJ�i#���TN�t����F4ك_kG-? 
5z�ؤ�KP>�SeF�6Q�[)�u�ʧw����mG��Yg؎P�3#GJs�Y��j�-�g	�~�r&m`"��8�NC�Ɓ5���~��m�l
����+V�#�Fӳ�3���g�!�[K©�X���c��?4�$�T�kK�n��Cc>8��k��S���m*!+�˿M=��iJz9r�$d�']�	�@n��7<|��#�?�^����9e�׀��죤�7���t~U����}��Cv�����d] *vW�DҠ�*����dM?[�(~6l��4Q|K��oF�L{�S|�_��Du/$��S�(=-��9aazB.�����J�e�wo�*�;��-���m�FLt�f6
O��b2*��!ۋx������>Q��EC������N����������?�B1��K�Y�]�&� �W6���K8��,�&�C��:�D�����%���>T��	�o�Dƻ�K� n�Y� �����M���b���e�B� 5p�*�$�W^\C���0����޺EeȲpW�!,`��Y]��s`iK5y��2U�TϽ&>�X�5B���V ������H@g{�7��֥u�7��d�Zy̯��5!z�;汛[؄����G�/��r'���\��-�mh�jP��d�p������;Y�����e�+#�JմC��؞~@��UHN�f2�P�j�ɪ�L~�|����Z:cE���0n�ep�&}Z봓TϪ B0�[�Q�v,�R)?���|�.�O֐`J/�!4!��򑛠(�(����3&��yLUT�E����&6������Աxa+�2c���&��sB��=KϚ�p�yPcu�I�Z$�`ᱝ�gVPq87����#	N)b���+�{4���2y��g��䴲_��:?6���S��ҥ�Ct1��o�����GR?V�.�|��{ʐt�Qe��&L�A3U�ޟ�{�z��}*���7�Yob�>��9���1|��[�Y4���j��y���QعWb�t|��(k#F��i:�f��(����2�df�W��n5�b-�C�H����}(���6�'����Q{��+Ģ�J�a��9˾}N�oh&<b 5�|w�+
��-�|���U�Q�- h��=�6o�3MQ�B*����L4l'NH��Eֵ�S1U-�S�-'%�H����r�U^��Q��m���c�⧘���{�e�(�*3�S����3����1<�g�ь�"��ۺ��r8n��}�����m˭����41�8���I��[�Q��I)����S7(�Iܢ���� :�#`��1�	��W3����Y�f�(A�����+�p�R�c~&�M�=P7�)�/��-]�mv{�n;�̫�54�d�NkF�����O�����z�Q=4#1�[T���8�m�Lg��]���/�Zc�'�����qf�V{z���g�H�G���ʭ����0+�a���'�����XF˳^��� :h��B hhdb�w�-A�����Һ��e�o�:?���J����?v�o���T�h�:b��F��&n+d�	O�)�)��+���f�Xk�jNd�t����
�P�s�,�d���=��X]Ɏ���H6Ѐ��@�s��@V�֎;>���)s�e��	��[-�=�@�73w��&���� ���?xp����P���O���94*�q���:Jǽ�!��d`��M@ /ۼ��7y{��h��O������f`+��/?A8����0t�;vp�Lf:��T<�|��~=d==?���n�Q��FFW��l>Ɨｊ%L����݃�s�Q���+�y.�-8�6��������4�o�&�Ό���e)�o�L�1�c�C
d1�X�@3�G�K�����|�5�)�κW�H���K������aL��Mf]�H�'dƼ������~ݐ!���O�(�L��hڼi֍ N��c�t���VF�Ձ��'9N�/&��R�n���1G�Kb(K>�~��Sg��:~?�r�!S����(�&�ŉ���*A+G���[��0;2���l�2@f�ZicJzB%S�]|x��R� �&K�%���j�>�k��� �pQu�U�0|a2�̥S����*�h3�`����^Ρ��%n����Ş�\vS�t:.��.����@�nW,@���X��TO��EV꜖�SՍ�`���ŀR�O���,�qM�F������	C��O`���sTp�J��Wd�c�̎1�h�XK���3�B��`U�����SU��Y��݋}Ͻ���b8IY�<��S�1A�� g� y�	�����Lٛ��B��q�7~���gy Wö�R�N�}=ɕ�ő��X���%���:G�x�W��	~������u>��+���x�%��2�{|��.�.Z��,���tV3l��X�Y��-1�i���:���{4�>:���HUϊFqg����a�1���m����{T~��2�H�D��&f���)B��n�u����: �Q'�u8�4���f���=�7f�ƛe
��}�e����x��Cza��V҅�QL/�%(� ���0Fj���QܞM���M�M�Uv��Q��h`�Zgu���C���,�	AgR���e��$��Њ��y�p8LxS�E�Y�\@U��N�s��M�;%�C~F�Զ���4�;��0�g'JJ.���b�9���u��|��o�(D:4\�b�]"�����o���N�9z=���e����Pa�r�w��Y�^��-#8:�<^Ӭc/���Q�o����z=U��v��K4l������/�ycq��
��*A�}l��̱
ҡ��.���"E���ò���h+�D�v$��)��2��vw�2������J�H.��=����2i%��U������j�Ur�a�T#��x5)�	�lY8��зׂ��op3�1�Ԍ�+D���@���t��*�CR�(�4��+[w�@�nQ;���;|&�$Y�N4'�� /;*k���,��o;hA��
m"z�[n��ռ��(�ei㍭^�N�E��fƕ�v��Gz~�ϟ����/'��a�1$�L��C(����/NRE����G��'�-#�����Pa��`��曅���긪'P�C�аJ	[Z���ė��㜵o����5�׏KV�^G�*Yv�I�<�+#е�#�QN�#1���֦]�H�����@Ƌ��9��<����}�>\���B ˮKc@� ^gO�tM-<t��H���$�d1��x�_������q�#���^�@�aL��`E��I��-Zy�s�q�ᓅ�p�>��� 
�|�m���F�u!&4;[�C�K�Z'�ԽO�ק؀nX���3e���#�/�QZ��y	�Vۡ���I>
���8K׉0��=e�h�_����T`�Z.�/�K�b��|�~'+F�@����D�єO_����*�i�:sc<�CP�K�UP�Qr̪rS=�����V#Uz�v�����w�ɀyW0"6��|!��Ef�K��n8G�j4A�lcw(Ēn�B�R!a��H����*�FQv�p�E��� ֖�3�%�G����N�4��Hô�_�?c}�� ������MXb�����C�����i�IFH� O��p�o�_ѫW�P�b�������DK1��n�T�9Kq�H��晑���:e�_̀ �/ґz+b�i�0�J}k��E�ܷ�o�^�>=�{��|�Q]�n���C�zY�ԋs�����t4ɝ�7��01o��zIr���Q�ѡ�\&梐Br� 	�(������9��E��F�o4�k� ��V�j�I�74.�s�G��&q�Yv�����~+)��.[����n�껍</*"�P�*p)���V��x�kl����43�S~�!8���CJq���4Cn��-����1Ҵ#���#��'~�u\� K���+��oM��z�~�g���j|����G'5�#�_F�p�4UD�=���v~��69��;\�e�8>}��t��8wb<m
��瓪_Wd��߹��9���[ip��?��$ ��qq�mYgR���Lx^����G�K�2O6�4ېp>~F��V�-�!fe���LU�i}�)����٨r��,R2���_q����sd�m��������
��K)�������,���M�Ts���-q��(#��F����Ɏ�2�ށ�/G0�3�OJ��	��]������z\�X�
>8˒�pT赮;�p	&���FoN��p���)�#3y�Ab������g��{�7��kփ�?�˺tq�B��C��B�^���f(9I|c�>��P��e�>%�QJ)��w�9��=||D@ih���P�7�l�	;�b�?�,h���J���S�:�\�S�X�[��A�cQ��Q����� �
��;|�c*���:��`�A���H�D����]۔�^-���p�D:]�|��X�/Ƀ����5a��Lb��^c��+8oT�7��I(?�PQ�������5nT�Z'��0������2�|R����vJ{d�$i4��Ġ�55���,��&.�g{�_j�~����FM �u�CQ�z/�GČ�-��	�Sb$х�bb%��ƚ��,�����)�.U�E�T�W��k��Ʉ�>��0�϶����@D��[�S�����������Ӏ	r]@9��*Q��lħ!7C[
7VǹB��u��ha��J�ę��h�ux��q���jAtnM_����$�J�U�}>l��N���'�p�Vy8N���S�j�`lG�!����l�H[�'i��G��lP����C�&["�fċ;��慈�%��EA�����:����L{�q"� j���e�JgyTM�+�\�4{����MW�e��5sE�3�0S������Mq�{�Ӌ�冟�c���6��*�(�㑟�,Ґ,ɴ.����6*L�}�R���_�;���w�������\�tU���"x�J*�}��x�\DP{��� G]�<�P�{i����I�ߤ�GvMf� �4�	)ܕ��۴u&#�Mg������N�pIhۖkL�E>"W!}�-vFc:Sy�&ceC��(y1Զ<qK��^�D��0���9�� ,��K%�f���n�
��>Z�����ᓅz��*�xA	���EO�-�ʡ�lA���b�j�T	��yr3��eOL�����S~�bY��-7>��"���� ��N��齩�LW��t�֤�{~�gQh�a�7�P�p$��"�&\�%B���沀9�DQ�}tb�g62�S�@8�D~�[xSp�:��ko�,!�_�b<Z�9��*{w ƴ��y�J����ҧT[�{۠f��IO�x�_� �!�ܧ.|<F�Þ�K�_h�?�YUw�����d�w�4\��K����4�s�3~lC�+y-��Zqr�(8�edn�����#�ƈ���Mc��1[i�ĩ��H�c?��踩e�Y�(���B���j˲����l����l��m�yQhހ��4O���7�a��h���$�#I�������, ����wre;�s���SkT{����������ȋ�%G���FOZ9������ڃ�|�gu1�o���υNĪ�.q�O$����nῗs>"	��pr�-Z�Lf���W50�RK���\_�y�D�䶉��4���}x{y�1Z��~5�`�4�+�۲�����%�G���X�5�v,�-�>���X��.>ޘvVd���¥ȯ�
����f�`��4�|���6D(뺞�a�̄�)]�Δ�~���:1�ݐ5���_@��;䂠�[򷺳�V��n��QjgX:�l:�@	��dc�W�U(bY����n�-�e�wM�P�dK�'���9yH?i��X�x��?��I���Β�a: _M�Jd��h�8����xN�$\�\O�/�Kg6��TV���dj$�EC'�:����z��F�T=OV�ɛB�5WtR:I����=5�T��@g���vW�7��xnGE��|lF/��T��t��B�1k�'��(m�W4�$��?�	��C��=I�� �CΛJ�	�*ܬE��V�t���9F�\���G�L�V��6�<;T�)m�yPͼ�b��V%�8eM�}��}U8e��7ɸ�7�m8gx���8=�>�n��MRVt�aN�3u���U2j�6�&���+wVG#���n�{	��=�^Q��q����˯�O�>d��wv���W�#��i8��MK���#�S�kT���,S�Q��sѽ���;�(����l�`�м�D���d�*����h,#kBci����EX�pT�*i�H�gu��fym��A�r�>��!U�����g���1>�l'���WzXi?7#���	g𓂡n��Dy�V���θ�@�^�?�2^�f_.N}~_��[N��b�F�`j|x��ϭ�(c=�Ӻ�ET��G,�R�*�M0�Z�p{� ��q�O�8p'���H�Y�0�`b8dX�1"$���Q5P��O1�%�}"d�g1����ᦒG�.�oj���l���Ն7g�*�7�{��+
;`���Gv�j[`����S��0���j�*SI4Ÿ�ݹ��B�d��R�}������0��e{��r�ɦ�~$ r^���&�z�m���A�
����g]���haC3�|!���~ɯ�#mv�>��Ϥ�~�����:N+>a���*�H=KWb*���v�
���b+���ф�t�Z�ڔ>|����>�����<�9+±=~�&�,��&��}��f^�_gj��쮑ogf�X#�<(k�f^b�G�id�#f����x>�i�FT,�D���������B�YV���1Fl1�M�����4�驨Nq�8�s�:��P�0Q���~�Z�Jv�8r�ݴ~Z!�#\Z�5�'%�(�9&�i<1��"tx ô+T�]I�6'�sK�Z�f�h�r�P�<���ϦާP'?�N��.hb���)xK�����_d|�Se�иq]��r+��X,�u�Uk]m˥X��*�U����9'���ߒ0���^ھ�d�X˶s�-��(˓V�\���A=z��W�D$���37t|T���-Z?����O�+����5�
�G�Z��B�7~q$9�'z��R+�VR1l��>�d���w�=c��H����q)�Y�}�#�fj��(���7�p�-#�Q� �:�C��#�9�,O�2�Hqa94kE��*#��>FΒ<x�`��šA$ A��ʍ�"�uB���ޅ����sƎ'������}[)�
�5���9�-�oج'��'�٫W����W�=��XO\VP��T�B@�c�GEhw<�U��`>��(g�R��K�㳥���(Y�`Ī��_��e:ۢ�d~EyD-OR.����A�4��^ L��s��}A��r�%�OK������d�V�gw�J*�_c!̧"Q������9����!8����
���6���3����׸۔-�ZӜ����F�o���dN �H�&�6��J�㽋������(�1�������lV����t��X��7;��i��Rd�ظ����:X�_���������?��+�Zl�$��pו^��_�b�ܝD
R)���)� k֜�-�AG��6]�_\`�WL� qvy��]p��>��K���J�AA[UwF %>0���������_h=D�B�j�ۅ6���,��Z�h.����:_�b+��%7���R�0?����f�y�����\l�W�uRNS�v�)\�h�%�kX�<H�m{�#�~���;�����E}�-
Z�]I����fH���g���#�E�o�4���e ��3��u��[�xV��t� O�E֮S�Mqf��F���Z:,�G�a��"�;Y�Ő�Il&�'�B�����xi�AW�%=��39�4˳�-Q���ò�����4��3��%�+u�+�J�Q�>>+���0�DK��
 p�e��T�]�v�������p��zRq����F ��9���c6-8������5�5J�c�� ��7�>�qM���ͳ�z�l���S �>ht%�8nc�{[9
0�q��� e�l�CeN�:\7Dt�)l/�Ҝ�5Y�(�V^$�G`�or��7M�@���yBRn{_T۱�E`K�qߠ��l������
)"K@2��a�]a�\�f{��6w'�U���U�0_
��K�����tE|1�N��!��z�r��Z��z7qoi�
^~W������W]^��<�d�� ��M L����mhDF�f�f�!���7���0
䋮՞d������?;M?�xb�m؃��=��T��njC$ ��	>�����t�i�>%�$���u\ZT��M12�u�l�������0�4ҩb �<�N��QClVv�Z��P��x��u}:�C=[D������w>�YX�8��rI�1߃�Y��|���Kb/�*h�Ej�s��h�"��RPS:v���2yE�dU���p5p�����`���-6/�<=}�
�L$�P%I���h�(8Fz�$m�����B^��ü���n󹫧�فp]P� b���>ơɍ���͕�lώQ�n*6,����NO��Ť�#�d2�oL�V����郪�7߁���GJU�q9޵����8A|ax;��~sZʍ}�u�^ՠ׮�X!"�0K��Ո��q��`Y-[���U{0�l�-�uFg��ۥT(�3:�»"��
v��Cy�_���D,��
h8`�ŶR������E��n}ڊf�ˬ���p=r��j��;2��W��H%)�7����Ok�.��g��KA�Pj>��.�P���B%z��0#Z����zzb����
�Ih�+�\�2;�/�����(�3*�F��DW�L�@�7&�R�"�R.�nkRs�3��)�S��%����$��'�o�)7 C��2s��K�3V��R*�n��,V?�M�t3�Q��������'������x�"���z�y� cH��Tx;40N�y
:/
�2o>qQ���{T��^%� � �=lp$�?��Ib��>K�Oԋ�EL?@�J��IΪ �Ƽ�?a�d�V�G(x�AH��pb+���Q���B<d<���4v't�$;�BIe˙��&g�C�����n)��zi�b�����TƜ����l���@�;��K�eK�l	��Rt��֗�]]F`w���5}���ؕ��Rb�?�ܳ�&�,��.Z�=��v�?JH�$+�vӮ���~���A;�L���οu�o����~��s�v�g�\�ꍧ*Y�ʵ��{�Ob>��?�m]�%94�B g�䈣%ʊٗ����iƖ�q)$ր���lOc�����'�����x����<a�#x���+�Ф�a�^&���/S*hۋ�!����hSG�^c�R�$m�1���E��ǔ��Y�TGr;�e"M���ߌ�˹ �.�ߐt_�B-����f���џ=����Xl��j���؉T�m�QD��o������1��ۓ��3`�E��X��Qd(Y�	vk��v���iRC�����\K���8�-�� �9EEL�\�E��l�-����Y��C��+i9O!	����2�&��'`�@'��D%��W�Ij��a��E�;m*�x�K��5ݔ�i)(��ʾҋ�d'��YTl'�C����S����,���E�w:��l%ᯀȷ�7���+=���!���X)�FO�Fjw��m-��s���KLAN�Ŧ�"��|����G^Ɓ(SQ�u��\� Z�հ�l2&���Ŗ���(=n�	E�{K�����ZO*���=H�q�Z%G=��i=M�q"�J��n�s��^Ɖ��T�Y�w���K��~�	\}0�H�ƍ;��<�.�1~���d
��v%)3] ����4_Q�qr��<�����u��e��MZ���#��B���*/�����5N�j��!I����N��z:.���pX��ЗT&>ޔ�K��g�W��~f"ċ}�!1��T�{��;�v;���-O��a���� Q:H�ҥ�y�ha�X/V��|���U�JK�RB��EQ:H��N �-[p[��>��89��F/�ް�rB$�L���c�H�		���/c��-q�ͽ�g�٭��*N�m����|�3��]Ai���U�\|��&Iڙb�	�b<#�?U@P]�>]�v{Y`� 3Uk:��p�k�V�AuT5��-O�Y<�(J���q����$��n�VoPzs�#����J��Du}V�a��i�E6�W}X�}����۽�v>�"(��W�I�P���B,^Ĥ�q��:����H���~�+Ԓ�l�뺒��A�nK�ϰv/=Xv�<
:�$ټ�8�L���Y�x��y�nM��<�zߺpv�dl8%���}��v%�BUu��g�v˘=���&�*5r��ؐ%���h	�8�,R�����_2zl���ic�C�oh}\p�1;I����l,BkI�xEUjN��#�T��f^Y�]��7G�˙�N�DS�)P���h+g_K���1}&��-���?��i�C���OMQ$�؂e�%8#=�^Љ������20%�3 �Q��	�#��N���lw!{���C����\$� oW��曕���	E��d�K(_�|��q~h�F[C���ɹ{��u2K�~�#3�@{7��/�U���O%GKG��g]��r�y�F~��rW�֎��Oً��k��g	�-�4����{�|��|.O���4�Þ��+��ʺ�.4�TJe��]C֛ɮ��i'$�	��V�e�������
aa��'�rH�����? uf��O'�$��E���("T��ΠB͛6�l][��p,�ݸ/ea���TTL�ܛtyQ�`�J�m=H�"m���z�m�n*�j�*���;$V��E�1B��VJ�]�# 啧��)1bN	��K�+N�xB��r+K���a��:�F}�����}=�W�BS��"n|(%u��>� �l?�{4��6�@��X�	�=%"�' ���#��"���Q���|��{��fvp����]q5���ݎ+F���3 9N��Y����n��jM$@��k���k�&�R�I���&>5�O� � �t���,A!pa�z��7���鉇��o�\���漇o���GY��pȒbvȬ&[Sw���G���J D�m�3���ѭ�۳�|{����7����@vں +⟥[�YZ�a�^��Ԡ` ��� ������(*�~�O�@���_?w�ǝ����0�hv���ήJ㜽C�'��y��S�a~��O{k�o�c�&O�����^:�5[��j�ݵ���@�G��&k|a��A�9�d�M.٭��b�PU!%���!}���Z�(�r��_�����Kmt:ԋbn�z�K�a�Y=�)W�E�pR��s�	]yyr
���A�Z�NOt�r��?)~O����[{3�,ٺRF5n���˩94���7�<�^�/~(�Jo�fK���Eu?g��$b�ҫ2���H�'�Jr�ۏ`�ʹ�TD��W,hkf5�m���'��W���F��F8�u��ǁ��D*�g����N茷�ޒVP�G/W`Ȁ�����C�Ɓ�Q�G�5�ɉ�:�":=Z<ь��_�9�'��/C�zk0�ԉ��WG��s�����x��ݗ(0�����%��xDuaU(���[*�Q�U���A��V$<n��?��uN�U�����8�9�6S�F�+����σs*�I���T� �
��v��u�`;<������IMTɌ�O=�+}��j���Vˌ,N�/.v��,K�S@2|�P�!�8߁n��@�qJuL7I��^jZA�z��袳;@�� ?X�&g�����΍u�"�!þwcaҦ�t(�� A��kFf��I_�̎���9	������&X�W�ƍj�H��G ���iE�
!�?���X��]�N!I߻��N��*֊L�����O���e�8����{am\Q^D�f�k�4q4�?{Mz�ab�����E����Oл}�gO ��!@Lџ�2Y�O�;TE��>z��Xz�V�N[��� .�/Ǿɠ)kMl��L|j�'(}��%���,�[�|���<H�n�~��nE|����"n��N�r��r��b�i����C�hu[�� \F/�}>�1du$[�����!�u����A_T���w�	
��n�Tb�Ek�e�wı>i��.-T^����lw@�wa@t��
�~���|J�HyU�R.+-g�k:�#�����N���LGu&eRa���li=З��J�9���A��)�W�-����¿����L�ߴ��6�މ;2�S����6���D~D�1��G�,���Xg��J�Ӎ�_6�/@I�������M2�S�؝�΢��~���0���B�dW��vrζ���ޣdy������<׻r�SP����-�H>��a/���-���h��R��{1�Ucp�BK���1zz�:��>��j5��Ʈ�;�k��ڐ�	��T�'����}�g�N�f���o_��e-�16*��_��b~.|���h���o��uf���I&$J
�K .< �j���tRQX�'���Y���_�P��a��CϤ�b��(�9�d�ׯ=tr�t�+���c��?)��󽡪-�
�[˼�ɟ�&:<��,���<Qu4�3�հu~Db�QZ3�&��vo����tzI�W��fߺ� �*�F&u϶7�V/u��1:V|\����=�J�� Y�ZO&�(>���8B��I����p
"���=�V`�pE�x�
����Kb�Q���:�9���i8�ю�����IګM�N	M�)X�먑f�!<)�$=�'���J����$���Gv2�;	�91�6�n��f
���+�ڳ��:�U0��
�1�������:7�ΏC/p��6�Pkgơ�(F�thw��\-H
GJ���9��Ńg���̕��Bc�|m3쌄K��-.�,����s[5��X��S�D�+�'��퉠���[a�(�w��>�K��ud�23�����8E��X}R��ҸV�1:�7 �Ђ��J��Z������۞{<?;h���Dm�"��sd+�d�m�kH��0pD3`�z�!,�P�r_ e�7�-�Q
3)D¢�92y\�il4�@�U�L�ؾ��9�;��F�HR+��o��@R�1XFQPj����!w����*lSM���q|@Ο���� H��_A��<'����b��×�� V��L�[�r�)x�EĆv�6&�Ǹ���>�98D@[|���K�_��hD�K���^2ni�p��{e���3�!Z�Y�e4FN�'�m�2v4:k����nFg,��+1��EA��l*f\d��^��Y�z�Đ
dz`O�(q�]O�-�Cu����Y'3_{���s $qa+3�l��W�Z�7ӛÖt¾uA���1*!ɍB ���Q�Z�
*�#j7��/����̴]��@��������x�E��c����\3k����ҙ��t?�E�oJ���fXhk�oj�/7|Lq�@6x�+%��r>ݙ�~��[S,��l)-�ɪ�uL�������N���v�k���#�s� ]:��_�p�����l��8/��e|�&�'�G��=$+�Ņ���R���>�%WaMV7;������X��4M�Q��DH(��Z�w�q[�-�W�����z��o>/QY���&[��w�n[�
����t�9�#����7S������J���cIQSlp2 4���,�oO�I��������Gƕ���e�"����L�e�½z^ɷ�ڑ9DG��d��e|d�R�B���G�g���˂hY����qS�Kl�)ѫ�yfZ��@?oܨ���0|�@���n8R�����ğ�i#�@�����q�D}q�������K-�IV���>Ɵzjs���+��>�h����z���DI��iO�R:���F�T�z��U��0��CI
���$�.K��yxm,Q^��>؜�p���_��m��_��E$HW�ϐŕ�M}
�5&�+<u$Sc�&?�"��*U<�@oY'P��k�B�'(���6´+����O�����;d�6yvJ�憒���Z����:�~�=�:���f0��񋆀��`�xZ��Alľ:��b�+�A��������@\���[�|��̌�-�vAy�uc����wR������L`�'�C�Ƕ��������0L�./�6��#���[�h,�晐p��i��4����K��6QRg~+�B
����݁�jd���L��t���z�S�%I�o�:9(�>=c�L+\���}�G�ܷ�g�u �}�P��xV�4Te�P1�F*�t"E���y��c�� �n�[m��s��֝���Тu?J��93�@)oX�ͫH	%��j�&���zx��h�^��ݬe��<��(Z�,M�Y�)�S�^���v��bi�6:�I��ى�!���CS��MrcRO����_�
#�`E��ظ�UP��f�f�o��Q�@��ǇuE���s����c�u2qf����&=�"f�OivF��E!XR�Cz����1��ar:θIe��� ���,�Tj��j��{�ɬ������C�:�C�m�$aW��2qgw۾hP&D�Wh'��nX���$���Q繷$���Ԍcjt'�@ߒh#��L.��X��]��,b��3���D#��<�/'��P���ۢlԞiS�+?�˲Q���g��{?	�Ѥ��*�d�`?2[ZN�Y>�z�D��TO���v��}���0�$v�V-k�v�pT�|�DU�|?!*�<�{ޘ%��y�O�Rs���)�O9 "/?�?Őt����ipvк|�)��@aE��,����6�uȒ��]�d�� �A7�?�%�=1����EΣ�={k�GA�J�(]q�m|
��`��4B'&}e�˥�h�
�\⠘RL�9IؑmT�4��7"�bu�Q�e*�>aްF��H ��<-ٙ�ҽ	�d�vޏ���A��*7a>VZ%�(��2'��XRy*Y��C�MKΧ\� ����@����V��Q��-A��:���I��7'��S�([�'Yt_]�y]=�n���c�C�A}�BT�I��X}����8��25'Z���H� ;��x_�d݇�aW�w���?���+���ۙO&as��~�5�s-0Me̊5k��p��!��@���>�-�C�Ykt:�+��A�m�b�Z�����0D7r�#���>D�['�|V�Nᎃ�$PE1�vtP���l�:v|-�_�iu$�2��z�/MC��Z@E0�⏾<���e)��+Z�D��P�~ز�<��<����ywX!�_��f� '~b+p�҃h;�+���E��R�E�>�
�r�MK�" �7p�/�H�hهX �TX��A%W�5!�$"EŃ"�l�l0-�lOp#��4g���s�c�����+!5�6�S�����oG�Q���6�����>���!����(�B��O��d�4GI=&A5���d��Ml��q}԰NM��7�'�S�e~��(APQ�<�j��s�.U8�����\]��2a�s��Cm�*��B&�Y2S��a���0�Ծ�)2�tJᇪ}m�Kd�8/ޢnXwX`� ��Qmpb���O����_cc�1��ӪK])��;0��~t#K��z��U�L8���@.��g�q틼)
��=z�]�n����#��/�|!;�H�O�ٝ�g�խ��
���BѤJM�Կ1�χ�$�J\�U{����h��y�-.5�\��q��>�a����j�	E�8���	�˛�b@%�g2�_hr�P��Ĭ��T���!�r^�f��[$4�ւ�N�SۑKu{��C�q;K���!�3
!p]�Kkr���G(��l����++Ma���$-��Jn����
��l�ѓXG&mWe�7��ouA��d5�S� �=���DmȘ?�˼Vo�?�^XY6�^X�U��?�s5�s���T�RN��e���^������X�Ef�K_q���)4��� cQ�l��Eke��T6<��1v���X%�q���/)M2+>π��a�{:�Z����?���B�C&�GDDg�۞	�ā��3o���o�;��I9�R�w]mK�@�P?��.s�H��c,����H|��[-��8�1��g��f�SN�=EP���Ø�1s���g�i�/����� �Ћ2��Y�x�	��+�' VA§L|犘¾n\�\����y�z��ʼq#�L�\��z��
~��j{p�lL}��ax��������1qJ?�o�`>"UN��+��ng	Be���X�HOu�R�q����v�CZߎ�/�Ց'l��N��7C��o���&�.29d�/j�>�:�­Z����bEY����@!g���ݐ�F��%�J�Ϸ\���9i�ܡ��KŬL��T���Y���Ϩ�H>�b��E6��-���~ځ�j-B�2� .Y�ϜSY���8P�TN��ꆂ�)4��[���������J-$V:<X�� �RA�̢ht�������M�Q5�$�����d*��~~`_	h����4����*��Kh�*��8�Ґo�}[&����j4f ��'	o�+�!�c�v�aШ6a�cM�0�s4U.��nS��⃨C\|-�c�L#Mh�_��$����3ٹ��C~�ԛD@@K��D�
j�3	?b��0x&��ɩ�ޒ�v�����s��ϧ��z�����Scfw�MߓT��ÎK��r{8���-���I>Z��=-��)�N"�lq"ZV�(�YZ��& G�'�|k!�\�d�h�U�V�`h;RV�?G���64�����ü�mV�ݭ�����d���%���m{=���N!�:3Q�x�`��K���a7��4�цԈ)PY�m��h\1�$�z���BXi��q�XU�Qs��$��*	�J�V�h�7���ݳ�g~��G.�c�ON�v��+r�ع#�k	uut�Sul�:�	@'g��^�U��'f��2���:�{�a+���ጆ����V�~�U��3w�<�F�R�rv�V`f��,�"��P��d�X�sļ��{�7bשL7Ol�.|&�Ks3:��������+�Cz�b2f�k>�2$����y�39m��`JPn�,�k�\ht�l��*m&��1~�e��� *�� Ya0�S��P��]�x�i�7o�~D]G���`׮�_�'r1��&�,"�B��4�:��9/W�]MQ�u]wW ��ET�xӸ����n���:z��e����TQ�Wz�a�V΋�qI-���.��[��,�X� �c�7���g~��0 }۲L�G���8�he�WV�!�B�5�r&�|X���/��gN��E�	3n�yn�&�d���~��%�XX��3���g�5���Qj�|mBu���H��SB��l}��K�yR/���y�ku~,�M,�89���5Z����&ɖU���h��*;��'�x�Țs�����NA�g�2���yj���F`�1D����O }�8��� Nj�D�����h�ϔz�Kd�+��U��شy&�|���-����@��9[������؊4Bm�������^/Άq�d�C��=�F`зq���K)�$T�.D��B8�
�� �����7f��,���?�2֐����C{��� ޫ������צG=�]����� ͣ��+�3z��X�(�u�x��+s!MIk٧�;�lV��4JQH`�s�Zs\l�**����Ǜ͇�����^�e�-e<�l9�iSr�+�%g�����+�M��#P�jő�����!U��-dׁdLO�nn�L.��F���dE!����}^"by��o�Je�UPo��lT��/T�)�#IK3�qwr�u�c�.�V���;5ۀϺr������A��\�eEA���nK��^]-�Xa2�\� Dem�w���K�q��fqK�V�pU5g�L��X��+UEЈuL��d\l�c A�7��1
^<\b��T`p�p��Ք�\�`�}��F�� �7sb`��*ܐ�r�ꔕ�& ��yBb�Ѓq���k������$	x�뢅v��,wqS�p��L|�(+o�#7ŗ���c~��D{Fhz7�[���@]i���t��2"���-�V#��H�C2��L�Ҥ�e�M�R+�������I���f�hK� 6~g���V3u�x�~��*�k�=���yJ��ө4��?�B2��0�-��&�	XwH�6�2�=q0�=�	��ه�?)��l�zmc��(�@|G�Kew�.�iʞ�-3�-d�LD�31���Z�2�-��gs�����\�e��i���5~PzG�zEyV北���\-�95:�J�c�a�~����豀�ΞMbk?����TG��!��R7��(������t�_H��_����pS�J�q���H���U[�H��^�4�L��NR�*:Hp(���)����w�"�+���;f,�sc�T+܇�H�x��o��fɮ��@��VG��Kg�B�7�v(l�g�b��Wf������+��%�i�8�:�Ș��7���O�hn�aU��*�0�%���R�vJ���e��;X:Q{a`���ܮ��]&��\�3]�d����F�V��NE��?s[���ł�Ox�a��C�l��<:Sw��]\gk�	4���P
�mg�)g��\FKԕ(8�A����7S#7��?����E�g9�ǜ� z8�N�r�����4,�����⇤�xZQ���P����_��f�\?�1�m��>q�����=�7�JEۡ�����B2}�Fi/D-�Q��=_�x�S0���b��)W%�>��K ì)�t2��+M�?����� [w�@H���	V���B����A�a�����d��xx�ṁ�Z-�?��H�ĉL�u<X�g��p~:��G};�W����0e����>� �`F19d����'8�+����[?�J�,�LEmx'�l|G�Cruxr�8N�4���HU���$E�)2y����V8���?*r^E�y�|� �J~�#<�C����N=���	o��/�-y��&�`8J�����@f�B�#�yn?2��c�9�g�N ϰ��9��b��o��b�����Qk������7�k��Z�p�C��G�3��_T���Y�t��*=؁�V�Yp|��mT��*��k佨p�-J��'�M����	�G��@U�xI}&ҽb�YIm�@PLY�/��f;�8(�2u����WkOEY��6��R�񖘗G��x�������A)���Hw��2@$��u��튘��Nrَ{CpN����N���7�C���u���6�E<�j;�Y%"�O	^�Ut,�x3tRHX�Ďp�@��R}��cu6���!,)��u?�u����x����"���ёѸڱ��~�{�h�9���*��/�Ж�Y���.	�I�EE:�b>5�RYf��OU!�(�_��á��)�2A��s��Kă�6 9B���E����o��� ���9�M����6ʷ�?�l(�m�K+IB��J���J'-r�Z���o��d��Ϧ����*C�f���S6�l��X��7$�G�B ߾M�8F�\D����p|&�Z�9jF�u�����/7���|;���{�JA~�m���
��������A�<b�9�y@L�A浻�1��!u��vor��d�sȤBo>��Z�����JHR'q����3��[�24F�&����(D]N�W��6՞��%q�s��G>X�=a$�l�DŠ�T�˧f�D�%����ۍ)|�� ׂM��ʍ���ṏ�x����I}w��6`>�y�S�po��Ջؤ�K�L�I��tK�H-��~�������9�HSC�V�;�t3��>o�S�F>����{� �5�Բ������P��euW찴�z��3�h�Nq,�史	2I_զ��"~�K�7p$d�e#��i�Ƨ�&5SX��m?6�P����K@e�;������AG�����5�7�/��/ �O�9�92j��%�2�lڛ�푨9��9�YV1�;Fʈ�5���y'��OR���iʃ���]i�L��/��Ws�ҟX���(t��7���fz4���� z�+�c�ߡ����8Ѷ]�i��n�<���w��H����� �P\���=џl���L�I~	���1���IC���ؘNw+A���96�Q�p��M�����,|�6�,M�_)d�V��Mb5oW���E�}���Y�Ph�"�\�3�y�X[���s:9t���\�Nʇ�w$�b��4��~�oZ�4�}!�}�]J����@��g�K��̐ ��!��� �ɐ<?Q�.��=&�T'��25v"�Q �޻SO��h�V̞E�(R�3ErҎA����K�f@��v�	��$x�)D_0�E\!�a�P5
{{�q�c��l�vG���c'f��AN��K	J5l:���jű(b4Z��=�)��(O\?��̎�i-Z�}�ʽ�h��.��l�HغA�"�����-�	g��bDI�U���͢΍�/,IU�=�q_��BW#�H(H��X|����"	��rPZ�z�`����8�x�*fR�_s�Z^,�te��,w�Fz �e'�f��
,�Ov��{�\�ڂm�P�MN�xjDwI�Ѡ��u5Q_	�e˥���� V�/m是�*���"�j�`���ks�uX�
�p��Q�c����Wԥ]�d[�N k���[~C��U�߈Y��>��T����|�j����|ӜBH%��ai�bvKv07FA�֞_U�#��~��k�9�Fv/b>p�������s��҉�&v�A�Q��:5V�Ȕj.��HY<V��9�zU�#���3�����Y�\?�Pax��`��� ���v"�˭v����@�N���L�y��u]������D0�E��7ݪ'R�ܚ=0 �H§���>�m�9�J��QyE��Z���ڀaL= �Y?s���Ҙ)����&�ĳ��%�4�h\gw�Kw-�щmuc�he�V#zc�c3���'BI1o�\i$uX���^�@�MP3Sf&�u��Z���^����w5���ڻ�{��� ��ڷ�W{�Ǳ�jC%Oz�s��*�i��R�ܦ�_�E��$�{fၞ\I%�M��E����3U��X�FA-Y0%H\׷�k��2˽:�u�w��1m���>4�e:.F�g��_�'��fM�E`9���ۿ��
��bY�I������8����,6V���/v�s�$@�*�Kt��5�S�~�4%˹h�!Z�n��:xW����ї8�hi�.��jM�����,,�4��,tن�i@r���@q���p��;�>=�h�zG`[�_�-`9c�3�sҬ⃕��^��2���$)*�F�Rһ�%H�;>�XEz��%�	
9�
X�5o�vx�:�E���I��58�ʰ�G4��8X~����Mg]��	�D��o2.2���j�q�|��!��dkx�v$]}x��G�&R�Ќ�T�g$ͭBs�τ �Ь�nw����`&*�L�]{|��*͖�FS�G�F{�I������S�U��cc]�^����!Jިo"��+�� �c���6s�Ci�?.�ŚaI���\��O��&X7\�l�X�4t��r��R��qx:�8p��4d+z��#����A�p�b��'�)�R���#a.�a�8-��9!"�_�1�$�1ؕ�Q��y��t�uh��ْ5&��F�,�r:q��|a���D��/Č��e"�7`�Rt�%Ż3"��N��Qz����a���?%o��ˋ6-,ƶ6�z�5=�!��:_����Ņ*�	�֙�����N�fΕ��C�I������K3n'+�3Se�W�%��<�����&�%e�䲽/�)�r������8w�g��p���W�r� ��8�r����Q_�y�~�$�foS�&)�l���44<�Y�8>{��?�n4�4�����#�
�P;�Zm�-�6��r5@�P���)o�h��7�Ex(�LVԴi݁�V����c�s�U�"芽X[�Cf����E��|g`Nc�5R�3�h�tS�C�V�eQ�7���W�B��M+e�9w:�����GiuL~���6��"��ѲV�_m�n�qVT��)�WS$����O)���aٓS=���Ŕh/� u����2������-x���R�ۅ<���ᓪ����۲�j���`�&_�ew�_���T�4^ﮔ����HXu����/���)z}Œ*�	u�F/E�ױ<k��neD(�Ɖ��8�)
�� �(��\�2�;�m�����s(l����m��_%m���v�\��}�֣�u�,$�e*A����l$b�n=�U�C�eCu(���ɔ�4&_������a%#=6�^W��t2�����k��쵓|��C�5�� _��G�h ��՘�i'�Ǭ~�~քJ �V��#���w���̀���`JGx/�io��Cwz����'	�h�z9.�B�_�b�ǀMɚ�6�o0=� vs��u2�+��$��3��O_=tT�����m��|�c>e$B|.'b4@���yҝ�;Z�.Z�<";Q�gh�Q�f������B^c�ء�C�Q-{�B���l�Ԓ�Uh�f��J��wF���H��+˼~ ��_�/c�q�y(���k����Yz���T�9�mp
l���N����*��t%��2�'g��@����Z��`5|�[�e%�I�Z�����ؐ�V�b�D8��3ټ���k�w�hx�ǻo�@nf�����94x� ���} H�3%;�m�*�t�<��:g�3�" ������@�4ͯ{��r U'�Y��Z�:��9k6�ѯr���Jb2����~�e���eR�CY�Q�/�d{��ü溿�~���Щ�cu�D�H��Z>��.� �&}�l�`��n��\­��l����:PYS�i�J�>�(��	����k�=(mX��$H��T���6.��X6�tD�%�3�� �8[�t����d"�x��i���[��OEt ��Gwp�7����عIf��V^6�-D}/ʅ�=��+�)N�[/���J���H�J.���5���]9�z=�1R�DsXc������˧�^H��TskRK�9��߭UY�8���e�1�D�X9�5绂zm��Y�o<7�(g�(��i�t�>a
YY����0���[O�;B���!��PO�i��l�e�{���A� '�8ͬm��	ά�eVTmo����w��:��J���lђ?�a�7w�a>��j<ĸ�I���e+7Jl�Vg&�G>1��ǚ��T�X�5���^�PT*��@Mw���r1�O�nD��8ƯQ K�2��ȥ��i�rH���JG��;����u��_��RaȅsV�I�����0��7�ӓ�@4��,��$ԝ�p߄Y�1�硂��V�%@)�>��������A��w%|�4E&�۲�2ё�T�۰��ѹG�.yX�W�PǉB�\S>��w2L�r�����o��ӗ�$��g�n3����0�ӂ��+g\$�mVa��OM`1���&��;�3���7�ͳw:�E�B��ڝ�р��fٝ1C��f@��VRp���m��o�H��L(�Dt?8c7sN����%c-�W}�����9 �x� �TdБ8^��[���T�j�� �N���j[]�M�����*�b�ֲ����p�`��aŵE���^��x�͘���-�T"Aܝ1��MT0�=�6q���IRf�yr�;/��T�F�_!�4|Xd����$f.���ٝ�B&�ME����hj� \��6��Z{!"K�gʩ�~�GG�T��E�hH����Q	�W��>#���U��؈��Rz�'�EF� �	����+�v�In�竞��;B�ٷ.�=b����R/|]�{��;��xg2f�pU'���~�K"����^�Z�$��옽V���N�?,ν�' �bD�Fh�y!�IIa��p#��eL�NBV����c�PO� �e��l�v٘#+>�k�Ps�Wv��U� ���K���O

ݬ?��au/:�#�oZ���%�����)M��j�Gb7�54��O$��S1o�3\�����z�uV�L��ΩԇƁ��FW)�7{k��V�Q >�;�k��P�G(���Dڀ�lho��& �l4�^�ߦ�H%�����V�v�%�O2B����#�fC�H�4�HҲ���<|��X� �&�([���~�?KDB�i+���2����X���0Mf�ƐA�Ƹ<���~84y�ZXbj DHǕ�wӖ��œ�]U�c�О^~g1����i1U� @�L���}^��#$d�3Q,��uF.E-)�d.����V���ͦ�2�e���+��ײ��.�dx���[ʘ(�չ�'T���L�쓭�w�����`���#nk��ҩ:ޔ�>���abK�gU�+ �퇒�q�H���0�֐�*�u['�j���g�DaT8m��B�ۗ��:T=��2H;v�Z��SP�[�B�k��|��!ԅʃ��]��>EL��ac�����'T1N;�E�#�F���-��=�-��aZ��n���	9�CK[&�!t��,���<���m{ޗ�V����zN���@-�xW��;��4���?�r�`���<��^A�NƜ"�}��,�2�weC��9���S
��=0�9���*���_���fOD�B	�X���v��l��t�[%X,��o����fH���=�Sc6m�[W1��E�˜Ѩvf�T� Y*�O�ۙ��D�PpY���Tlԥ�D��-]{z��s�5���~O� ��U���fC9l�X4x^{ʽ"fN1�L@��LA���w���ݺ#�s)C�K
�~;��?�!QC�GѨ`?��c��o�*_��P���׹D�OU)�č�.�������@T?��H_�}���s����S�����U���b/��[��ί)�PFC,C1Ƣ��MrS��;T��'��QRK�]�����Rh/�6���w:_%Ҹ#Jq�J�CNO���vhk\QsD�mֽx�N)�>}ι7c��Y�e�D�����7�C��G�$@�A�m���XB۩ᓾ*2�ԴN�JK/x�;��7��B�%��A��h|��0܃E���$!'U4Ev��t�����Z��M�?���%3�H�5����.���ŏ�߀��9���oE�jH��C�+"��6{�p��T*-����3�V*F��l��&	�^��H���A�E?�op�!���-�0%p
ص1�ڦ#��n�=�[G�F߿�b��~=F��W��w��Ԯ�dCtz]@(�%F?���%����E����}�}�s�%�0 �/�҆�^*Ω\q�=:0=�d��u�[]�K�j�1���EԿ�pB�����o�h�S i�N��Ǿ1��2��&���6�Sj�9����/�S��0��pS�q���}n�55�QK���KDI�z���܁F��k��<�y�إ5ԫ�l�}�{!��3�������	�)�����	������tR�y�+fxW�&<O��Ћ�x��Y�;���ે���-]�@<�qT{���J�|��o�ҕ�m��-5%Bǵ�G��uw�}�َvhpqنe��ڄ�$d�p�<|9y�fI�yXL�;#ߍ���̴\�+ܷ���pM�!΍P�՜��L̒6��y��i���ׯ�D�M�RӼ���i���]"�FI��,�����]mK�৅;��!�eMY{t,���r�
�a���5�Y�E����	�\1n¥�*#g�Cn�W�*�%���2Dph����.���oFc�`��@���ߵ[�rԠ���0�>���a�&��H���*q.�:���^�4)R��܌���qF����i�׶���n7�� �K�C�X�>!���\B?�'����9�;���Ƌ��0��`��=,�t�.�\�v��d�������<GϡW��������w����.�W��Z@UmD�<Y6��Ԛڛz8T��i�'�f�{���}+�Ԯaܘ�^G5��S��E$�LiT��b׈;���\j�`�?�*�u�=�M.��N9ˋ��W�LP����q��xD�ڬ!:�z 
%�����qՅ�ؽ8hu-�>���h�˂Ip��y�.�z��;eI�����;`w%G¸���������z��24��3��ܴ}<�� V�|ʑ�F�$�����(D���
�0��k,ǀ�F�o��A�����` U�`>L�-Q�*�)Sfy0C��X�������M <
�F9��.��U�js��^1��:����2N�sc#�&'��b5�/z���A�R�5#kkH��g4
TK�lP]�k_��:Ҡy�ߒ�������a�d{�5�����Y'�$jM�ğ MӴ�J�6�r�GV�$�b� cA�T96�p�O��:W�����TXc$W �
O����vD#��Ѻ6�z#�$ =WF�'-�6|:��R��jd�{^�A�ѻ7j�jpw��R�y
�4��ꇳ�02�Ω���[���9	H^*�hW���p%wЙ�-���*����z��ǁ��z� *\�o�N�!,�����)nt�5�`ڭ�5J��
ɺ0�2������zS\��9-b��N�v�%< ��i;{|�QZ ��K*����XE�l���\Ⱥ��
[d��LL�S�l�� @���?lX���,�h�7gQI�&�r��I��_{�k0p�7E�߰k���hG]�[э!����G?���4&�d�,��1�D��N�/O��c�O��}#?Ι r���4
J9Lj�*⪊L����˽#�6��gk�$
���A���Ѳ����]%){�_U����)h��]7���7���Dje u_w'�E5g���p��&�%���k�N��!�z�C�
R2wq�%kē��`�@����W��T�$p@�}><�d��흃�x�kԟ�	���:��::�wҚAz�6�{,�&��ɶ��F��(��Te����;�I�H>~xP�n���B����J��,��4H}&S��]��!P��kz�85m��%���u�!��>N�H����'g��d�dƖ��-+�y9�8s�<�i���ؔ���P?�����	�x?���r��%`��=d��B&{����J�T�`'&Y��]~*��J�؏�wU�@�IZШ�%����9X���5Ȉ
�d��7��@G΍�������1�D�a�y���mTP��J�o����+"�T,{t�{P+,�7���ph��1ݐ�F��\%�*u �������k�'�D3�����f��-QX��G|�qC�ƌ�o��Ju���в��*������q�Ly^
�6��T���0�H��?��'�̉��B��)w��u� ��W[m��ؐ).�M��I������ ��Z�Ԕ�?l�(�c��v��	t�P��jOq��^�̟�C`��fr��R�`Q}C&�$Pfo�����".�p��_�9*�m��R�}�8�� &M�����햦��2��6�|q����F�`Ä���lS�,�D@I�W����t�c�#�)���&�E_�zEE�bAqh��m���d/�$� ݒ�O�>w�Wy�� t���"���`�C��Y���.�9�إ攛ҰyX���������|Z���@z%vo�@�:���w�<�LO����\�?��B��RĈ����n�?�5�E0���B!\B���YKf�Մ�po	�0��g���W.�Z���-�x���,
�d�]��p� N�� p�U�)�2A��d��#y�.��nZ���m��0��.ZF�ݫӸZ ���?/��A���n���>�~݁tp�1b�5�����c��	�V��j7�~�mn�'y1��{��K;�]�r�-�Wq�N�g��d�{'�<2w_M��*�9A|�_� ����
�s2K��W-�\$VF{�,ް5�",YU·r�N��q(�@�������X�ӊ��N�����e`����9��Ҳ#��x���nP�E�.=�}��`�Zx��*��8t_�z����G}���_���	/�N�G�o�	?��)�b�f88���i���zO�u�9���`�z��� ���!I��Q9�Z�<���`�#���?���Wɲ|�p�@G�4nYjGy�o��ڤa��"/r�б��A	�i�>u��%7�'(a������I]�y����yi9�roa�m>k��:�\��w6���>v��nkկ}ϴ��a�K���X%˺J�J��)[
�å$Fd��-$��3�����f�Y���$[��c�u��Z�M���M��!���x	՛�����e)_�O�B���ac��LpC%���d�ٷ#Bo��v���T�;&����&ڏ�VG2��b,Vؙ�*B�\ƚv��}u��e
�t`f�T=\� F(��i, ����`����^�o_�>�u�*�yP�2I�rZ��i�đ��cyǁߴk�����w{�g;���j�홃ʊQ_	����l��R��)
�!�JHmSӎ�[p�i~�n~:i�r�\-�b̵o�v���}�E9�VY���ܳo��y�)n�G�ԣ%�`�%Dd��yS��A	��b%!"U��;Y\�C�5��'� �� �����
���c�q���w(P�z8N"�2dpV���=$e`�])���H�l���6�"z���x��M����7�c�x�Ը�����(VUq�V�!����gS�z����9�N	CiL$�i��U=�U��>/����q	ܰ�ɮVIᬯ�r���B�O���E�~��"���%��D<�wS�6S�ۂ;����p��!�����/�-����T��1A���1{��&��}��$%��E?n΁Ŝ,��2���
Sc�DF���pF���,��o�OE��,���p����Ê�X�=P�њ����5څ�ړ�z�j"��4�L�QB��"])YK�O�{���"o�'Z��Ѱ��)�5������"_!=��~G���蠲)��-&X �������	jr4"g���/U�`����7�g�.8�M2�.�Ɍ0^����i?��*U�bPcG��"8�h��K�˰�DS`�g3�\z��2[zg��� �׽>�� ��n��K����w?e���MՋ��b���e�p�3WW� ��#�W�P�PN@i���;+3��e���|��tՍ�z���B�)�HW Q
,�n&�n�Ӥ�qrܸ����� ^��>46�Z���s�.Z�D{�1�������S3ȕ���J�)���ԝ���4�eҧo&L[������k�~V���j��K��%/��@-��=��َ��EG9�V�=$59)r>���Kv(A��ز�-��9���D�.[�%m�! �i��,�ZW��������z���8吺�c٥6CE�ɇ.稺��%S��?���k��q:�Ԣp.��W0�vPʲ��+�r\��yJ���u�7����o99a��vm��8��l� :˓���y�{����y��W�cN�I"�O���/�t��&�{���3I�/�8�F�z�\���L�`���'��s��D��o�EFY/Οe�4�ҙ��B�8�h�OE�L��E���s�ޒ6b�I6>	��Ӌ�Ӣ&W<2���2��p��
������!���U�*+'e��㡴#�9n�9M��M�[� N�C�ݬ�q�p��7j���	�����2s�>ݑ�475^��6'Y�e�3�w�-&Y�L�G��XFg_-�4�<ދ�K�;�<���RP"�I���^%iv+��ޜt%B�g�,�U�f�J|O ���tΫ���n+Ӫ]����Ѫ;����M�	}���
˟�SU_%��2��ђ�ҫ���
,uGG�Q_vW�"Nꍕ熂y/���'�9ȫTf�6 ��r�x�z�\����?K�W;���F�p��$��� usp�Ý\��`h}?2��#:���<)��}��q�6��╨�����������6"�@-+;����I��p�[n��SNV��KPo�DQs��&6�3�KV�d9���h\��+�c"���>�@��(�}q�(�i�m'e�֝Mii���!��bsv��_kC��8,�uo(tRv�t�>Pk��PSv-X8�Hk��r����?B�}B�°jE<�o`X��PG7�X�>�� �����!(mm%�£:(>�
�d";�gF'�h�8~���sHGt��[C��|�1��L5�c������)S�l_^,(钿n�!�v���r����$�T�q�9��8�"RjH��C���$�]0���B�si����9�Ǩ�gG-ҿ�ӌv# +1�-lN �f��:bɶE�~q��2���r��FG���8�e���wGLn*n(R����"�0ͭA�h��;�Wuo�Śi��U��I8���67�F�dC��,���Vs�A'�w�)�nc��+؊/�+���\N1�6�,> �B�a�"��ya&��,����h����9&��Qƥ��c7��|�ՁH��b�j��aȒt/�TO��0,A�ǎ	H>�;��x���i��7�I?�gv���N�E�h�[�ǽ�̠ֵK�ۚ�D7s'�����j��� ���l�����7N܏<�DK@J#V��J�QCNmh�4�x��W�u��[Љ��>�%�Jh��ŕ��#;�Q>��aj H�[QI�#�͗k��)Z�=�˓�H�RG�1Cֻ	���Tg������ҵ�,HQ����Nt'�b3CI�b�]���i���rn�G�K�PTVK��v�؛�ns^Q�&����0���S��b^������W�Q�ha��3H��T5wg�ʱ�kI����1�49m�C���+�x�����9�1��r�Ngd�?
_1�d"\g7�3~�!�ѷ�f��򮝬=K�j=��e�;+��k*�/��U!�F��O��U�ֶJ�ѿD�_(~b	�r�g��Ns��z)?��1>�KxU�Дs�5M@}�4���W����=$����@� @�n~}�^� AG�4��.��X��gk�&-�/Ե΍�'��f��7��~Am�����m����>Qq�S���@��E���Г �cEQN�[s�()	�A5?��y�9��tb";�V���6�RJH��
�*�+zd4B�xЏ�R%R��6D�÷R��"����/��l%Y�g��Mr�����ʶhF�X ��o�ϙ�ee���K��nE:���k�#�dۜź�w�>�s��r�^�a����X�û�PQ��g2"��A�Ь���C� ��{�_�J�Az�#^�V=⣥`V��0�sѳ���Q�q��q$��p)GR�����(�-�{�3��T��g��G�����D�}���l��ahi�hL����o&�#h�S�K����(*'D���,�=��!�	׵/��r L&�>�O6��M[#�߬-h�3��)1�)�`����\�$�u��ޟ}>LdI�}���c�!��W�� �%1nm�������|�E�I�l�	�62����NRݲo�2�J�W���)���6��ۜ����&���#�m�9�?��B��ٕ���Y=g\��,l�5��&{��A�F�)���X:�t��Ǯ=���0��D�y�3��\:��XV�l�����o:�`V�jJ�W���k���"�u����ݼ��-���L"![6��p�L@2�bQ��d�|>�pI����TD͋�rE��L�`?�}?��:7��MA�v���IUH��l��.Y䡄E�
�S�g�5t�,>�*~~�p��M�,����WC��L��N��g��,�/}/>|b�Sj�pU��P��6�Nq�ǞǨ��-��q~�)�����906I�c�D�)�[�r�gU6����C�x��Ri>���rsJ#]��';MS����J�����4��$���C��_�*CD�f�&з� BF/X)����mOf����?yb[��w{
�!�C����k��|[(h�8�������:�'�+��0l���U؛�2���rOh�l[�\�c~&�������`m�2.���E����v���χ�+���%�Y��ce,� �;A������� ޷o.�g��*�ɳ��VulY��b�Qbyn`n��Ш� $��}5R�/kL���\��}_|O}�-t)%��^7��X� �Yw�^1�i[��?=<�j���{=X�9�����@r�L	�CW���n��cI�J�I#��Ҍ�d���4�GNi@Iv�����C��Q|B��a�ww�W.x�@�>��
}�pp��	t;���7/Z���Þ�o���&�j
�ޓ��FS������n
�h~OYf:�$9�`�\V�}޷8˒�_@�5����[�O6������iJ��9�� �@Ap~���N,`@�\2�\�j�0��"?��J7E�lM�2��Jr�7��ZA�������*�^�:)c�Ǩ����W�eb�^T��6�x��>��om��;�Ы�5��%q'`/�?�xBFk�2m���7�*`S:?��e&@�{#Hz����6
\�y�	j,�
���~Kl@��H�]�V����Mt1�mY�G+�B]�l��Z��ب����m���ї���ug�2�;�mt+h�J���/r�\����h���evYA��PRd���S�:5��m��[�1��K�
Dkzj%�ػ����;�T�h'��-VQ�g_�<���.�K�1�u�s�Y��=�d;)������
B�0��K;�i��<kQ�i�W=U���v�11jU��,X���zB �w�F��Nru��j ��R���ӆ�i7�(Ir��3s�2ʧV
w���-�ѷx�j��㚦#gh�F �tWć9a��~�ާ��e�,�o�W�$��n£��K�Y"d�}"���f�Y�?�ጌ,�ڴ�H�*�s;���c�#��X�^$՚-�s���+��2��ʜ���c�B.�{��($��f�-rpԗ���(x{��}ˇ�:Ü76����M}i�2�������Þ��JC,��Β��eie���܁Ŷ	�n�J[�U��K]se��'M"����'7�@ɮ,8��P���yb��"��[`�з��q�i	\�gp�cpe���M~e�x�+:e�g4�uH7S���yxu]��+�G����^&<�6��ϩж��F�pw�\>���,����:�0D�]v�Hn���J{��f\�qp�װO�z�R������O��?��g�?�2G�.:���������{�올�M�)s���1��������k�S�н�Z:�r�(�|j��w���n{_�z�M��4�"���B�l`OiMVV%$���� ��4���n���A7,��A�e׋A'##ũ��RGs��������e�Lb�
�I�\�ڊs���ʌ��:Vյ9�Z�ȴh�0��у�'w(�̼��I�α�mW�Q�v��:�Ѩ��c^/���B���?�4놏n�I��A>��u@̌n���i��{�ʎ������@���FN+ΚU���z�MŦ�A��aӥ�=A�6�}��p~���R�O��)q��^��������z��IL��s�$c���U��%�J_}zTv���P.�J�fV����6g�D�D�@/�Wα�~�/ֽ'h�>=V�W�s���#��|
��˚~��K�LM���3�i�VE�.=9c[n'f�b�~1!k�J�h+��'�4�wơg����R|>���4O�2��L��iS��^�1������B����S&��?�{�Ѓn몋�X3�m��cRv���a�H��o#�Wu�- ;M���Əb�m'v�]I	=��z� �)}��ᯨO�|av?�~1%}�����BGe�ai�I�Ǯ/��F\��?�`��~��.��|d�6�<����9�e�Kqyp�c�ͩ��X��r�(@��5��K�����Mܲh���|˵ȵSҪN��i�bؖ!����#�l�A^���8+��Œ���OH|o��ĉ��=T_�W/퀴��]1�V�؈�?����T-��N�I�dJ������[�)���Q�Tۧ����.�E�*���Ζv��jL�y�KS;@�M� �f۽�V�<��)�ck�d�F���0��|�-!%�n�Jr>te�G��ӏ��>���pqMʧ<�z`ţ�qQ�Leb�W}�lċ�,M7��Z8n��C;�<;X����KD���2rj5>-u���$����2"ǹ-[;��;+���j�*; �W���u��>7�a ]ܛ���c�.o����N>X�	9�5�4u�a?��P���ȰY�h����c����S���e>����
�h�����`�G�����)�wV���yi����s�&�>�<W<��p�kb��v�4`W��x|�k�g@�h���.*�έj�{�SXK�G�$�JF�
��?_��3�Q��}.#�ܦ%/a��S�s=��n����Y�W�þ?+���Ǽ@,�t�)��|�������ֽP��F��,g��S���J�ʻ���?'�y��Ɨ�DW6�ly���Iȇ�	8LF�e���0����#p���Cr��݄=�1K.1�����Ӡg'�P/�P�)���)ֿ2�ZE�1�Cg����W+;s #V �&�p�m-
6�
��b���T`ګ#�,�9���[x��˼�E-n%Z�i�1�`G��.��eF���@�N�ɟ��Hs��*�bI>,��r��Ō�	6���s����2�G��霈A��i�wƷ?����Ow˒�����v*x=�]Q�/^,{�5,Q�(�z7L�0f�E;�F��Cޜ�`m��h�L�bf�y3h���y
�	���i1V��Z	���*jh���a9�DAs���E*Z�����ևY���U�B���u1+D�ڐX)ʓ���)F���=�����l��I����1 �l`a�d�B>��P�:(E������T�bq�&]�ΧC�jӮ�ta�-?7(!�W(�z������#w��ĵ�Ӥ��ixx����EL@ܑ���2�t��
6j�������ŤP��_=�f,*�H�{zĖ>��y�(��4�;��M�i���?<�MQbrE;z�.�E��r����a;ĖopF`Pbk��%�����jZkS��F���QrE�C!�
�]�f��?�����>��d�a8�i�bGdQK'CFs��T���G�|/9���R�EJ�H���ٱc��s>A��6+��Е�6��ey��3���� �R#(I0+���'�����F�h��u��͌�Es�N�F=���@�� �QL��t���pY�=�V���(ꈲ@��6����0�a��'Tq��O���
K�������m*���-f�0
�Co�����y�f�rdY�q�G�V�Y��9�2�͟���01�I� ���-�x���L���/8;^�CBT��E���n�rcs��!�]DFul�yW	�8�Kp-��X�V.��~����C���gL�r��!�	�q��0à�r��Z���h��."���k@���Vj�1<!d� ��K���@��ζ��qh#�E��h[M���Ǎ��W�j 2��!>������j��\�j��|��A�3���r`��/��ts_��|rT�o	{�q93�l�H� O�dBf@������!����E��*l��s�;=ў��)�eF���4�$xj>%�,!��|m�0�J5f;O�kHҌ����np���6�i�f��>y�v`��ȴ���R�p��U��� �������#5m	��S2�0�>p6x��Xlkv�A�o9�� ��Wd	�mq,�8܆����C��I�D�b����{\���ibi}ȣ�D�b�8Z���e�f�}Ea��g�7M�����"��d�?��d'Y����#=T��ya����eQF�T��y���*J	:l���b�Y�Ȱkx�[��Uxŕq���&![�OL ����
������3H������l(�,�J1�B}*mb�;�h$���4Y���D������{��\���0�f��*�����AY�l�jT�� kN���D�)A�������S��:��ņ�{��[06��c��VbNߨ���5���nb�cዚ���V��b�����Yw(�ش7�q/���7�I}ܟ��3����5�Fz� U�km�G���ºa�x�u?�l4:� ��XR޳��M
i"�J��c�aF�y;0zm4d/H~����">���6����N\�C*�(�tV��p��{�;ym;�+.����b�h��m?�<��l>[�F\��4>��&�	t�Ps!����Jе,�/�w���0��0V`��?mgj��0���L��!�N�P.�����S��k�9y6Y;ԖR��w������r(��KA��gdt���L��vIB�bY��0����[�����վ�j��'����<�YV�C-}SZI_ D
�����9�,w�0^��g �ވ�����̶�J&��칓��Y��{1y'�p��.\/�g?Ã��޵�\n<ܽ������28XH�+	1U�Ѯ��6"��r�:e	��a�!B��*"b��3%���K ��\hݟ��c�7�g�@G�Lm�-�/�>�g�[�
��+�Ƽ��O��M]Mߦ6�v\䛥ήW��M��[���y�,�k(6�1N�TQ�ݑ�B�Q�wO~�}	p�Ƅ�E����D�]�9/-uf�o�HCE�CVU6y>QP�-�g���_f�c��X��8v�Δp� ��#(?
B�}�ل�8�@�m<���ݷ��.���_d��cΔ�ok�d6��WVLzd3�TZ�fT�$�b�+PU*��;l�.fs��!l�L��%*I������\����j��E���f��0zH�
��ڒe�i�
��v�`����{�$h�0��J!��B�B� E�Oe6���& ���(��0$�Lk���z�b3�L��l-�lB��K4o�c��׮��I���7e�6����(gI�T�ٞM�)�Zo�q@1��^��WU����6�����P&�X��ٯ8�nf��$C�g��+�	�O�����S�K�+�
!u��!i�I��aX�ƬR�4���O^� c]��U����v�JT�^��d	0���2|^[�9 �����0��X�V�*�5��>aC˭�q��}9��ƺu_�bX��lE^�R��I�MB�w��_�����#���[r�j��	�����!�g�-��:%��W�
@'4?<�Z�9*[v��"�+"����܈-{h3�1�l@�Ձ���uDug|9&��ׁ�&���e8��ط���2�B�_v>����W̌����Gy��4��R-�pd�g]�;J���s	@�����	� R��b_1�|R�,�i�Ҷ9ݖm�)ë�)bn񟶬a��z���z"z�8r"��f�гE_�ڣL�m^�,axKX���VT}��e���WJ	�QDo�Wk��|G��6[ݺ=�c����H�#Ʃ��wH�s�@=�4��$,�
�?S�E���h=�[l�Dʋ��>s޷��� ��Ib]�3�(�O�U'��ߑ7��~��GZ�b�!+E52;�sGx��+�Wb=�c��=�Cmd�}ù�SW`Ȟ�͉w�g�i>�&V�Jy��1Mi���r��L���S�'�]�ܟ�+�B�=��ñX�HO�@dK�|���"�:~X����X��( �s*�Ui��!��,��Q�
P/0�RA7a�Θ��<��o���Hb���*>��v���~�m`O��{�Z���8.Зe0B�?ɡ��XȠX��K��WKG1�R�|4Rzp��Ȃ����)�
��,wz�����z�ّ�\?�X�{���ք����k��_�9=��D���\ݔ��]�����_�vk@�eb�fޣ=�7��i�S͞M�`QŠ3��X�GO�Z��4�� +��-�7���CEv�����;ܰ3��`B���>1Z��ߍ�y���:��+(B��N��W�\�)�.�3�P�Gw�*������
@U�IM_,�:�9�D�G��OU#�8B�l?�� 6$�^�n9��+�׮�U��]��7�2�c �+���yO\������|���'�JK�����fL�t5]�f�>[����c�q�d�5A�dX00K[a�:>�IBw��:�2�� ����,��t:�P�gs��d(�V���b'h��m���G0Fj�m5{ ü�-����˓�����ZB֐��v8હ:���e�����#ܻW?�;)m}dtH�+/�J�f	VJ�J�b�W�����=Ǹ+N��IQ���E"�%撦�$�͞����H&L���0��*@���8Ƅ�)G�<�K���&'��Q*ps^H���	�b1X 6�y��~����+�
p���?[�&w�ِ2Д<�A8Q�Es��H1"��V��Zp\p��:��l[����'ՠ������R��w�Q�(�S���W]û�kƂ�v��R�cc��jd�Zp�j|<���Ĺ��jɢ�4��1v��(7U�/M�#r�Ȝ�hY��� �$��i��c�
C0�tH% �Ďxbt���"��Z~� �&��N���%z����9�͌�,#F|�r��r;o��v�~�����F ��64([g���y��	&��P�m��@yA�����R(g��a�܂8+����c�7s1�P�XQ�so�Ro1�|s,�6֒f��T6�`�C;��vv~��Gq�K��S�]�h��a��d�8�nRH9������W8bH�U� R�Y!E����s�&1��#�h�'t�&�ZG��h�X�yB{�_�צAC���\�`�����v��}Z�Ǝ�H	)�E�SK*譞�D�I�ޤ��g�:ǟP�;���ˮ�<����Y���{ݪm"�:�K�Ej����!w�@i��>�z��p��*��P��#���>M��Gi'�[�9Q��^�:�9�|5,�o[yi|��Ȫ�T��&����:�����a<h��Q꾝!
�ۡ~хV�KP��Eg������3����V~�2��;ū����ERW�c8�wp�z�!���ʏ֢#��މ��Mv�S���W�I�����#.���
��o�M/a���_������`�W�o����"��Ey	`:�S��z	{�������ӏ�H��nzi-ӧSw[��W�_�Y��M���<����bY��D�w�L:�ă�K*��j�Ei(��CO�V�t�^i)N�"�;����e�kW^����y���YOA���	�+0���Ӏ{/�[�x���̽T2�9�56� 9��%r�gǏ����w���\��s�'�&�:�b�n�(�*Zx��z@ҲPl�����!\��XPD)M�����v��s������pj�,vK�AT�Hdx���*sZ�	@(|u��I����Bp@9ߖ:4`�%��c ���Y|
�<�� �%� "n5c2M�!��m�19)���a7C<��������GK���A�Oz�.�k��:���~�Q�e�fO՜�I�͒Jc�+@��[_)��l�t�S���4�l��w�M��͈/J�&��3k�7��(���<�y�a�<�V΄n��,�Iၞj��j'D�U�4�����;6�V�EW���q	W|�*6��	��Ԧu.!�Ҳ����p��?���>lW������§��w�3
i��s���g�s�w����3���a�x�UD�ʇ.�,���L����!%Y
��KF~������Gkȯ�n 	�*�T1j/�p��L7�@F
�O�I��F����@R�{{nYZ�H&��$-|Y9�/9����U�M�^�,�h�~}:u}L��0m�H�V�y+��pg����HB��*�"�֩ʏh��8�
�/�aз�G4�U��'�D�|���i1�Rt�R/gEK>L���G�IcI��bl�P�� �WC�bg�F��OP�s��~A��s�n֓J�SK�x�)ր?����� v\�B�Q�Z�'�;�E_�i�p��`^^����-�!r9�u���e2=���5�qU��D���K&�9�!%:� Ϊf6a�f��a�ĥC�+���!�{�[��a�$+�:d��=Qh�z(+}��k��
34c���L�=�����w�N_�@3?+��[/��5�'�����9���F|�I��
}x{��9��pF�O����#�˱cb�B@"���1���{B��O!۞�ݥ���%�#���:*���I�9�s�ތ�(4�A��F�������Қ��W�]��Lj��Y�@��a����-�4�^?b%�����Ѓh-eYA��@�\�������P���p�X��_hq&86�0�9"�G�|$�7��B���f.�HR���"���Z*���!�S���#V��<b��O�#�ǭ���'���J/{pE������1e���D�dӅ�m�[�)K$�����W(�2T1W���9�U��]�:��ޱa7f��^x�D]�8�6\G���V�FQX(xK	����׀�$��K&��m�M�I
���:D�.BQNP�$}T*W��.�����˕_O���~��v `Q�W������4}&�)��;��[]57o�Ye���%� ,t8/zo�#�_,�@ev�s-|�� �s��bto��4̨�s*�n���n�FsjV�b������� Z���g��M�rLZ���Tp�F��*B���g6��}�U7�N�>ѩM�o��H!^[�`�
��
h|���P����x�l�0S��ً�cz��5
M|���̖X|U\+}3���f�݂O�-������� *#f�98�!����sU����\�B�(%r:�1S����3*Y��RNZ ��Ǥ�>U�T������]��4X��(�
[M㲾�8}A���!�٘=:�m�䤽�	�Fg�M:���`TX�t�o�$�&�����q�D�JV/�X��T�U����۠�����D0��֚�[�:�a�$�"���{�=�I�d��X�I�9�ȑZ��Bdv�.? �ٵ��hݒ�*�*�!3Ӵ-�0k�v$���\�:r�ϥn�ӗ�٠M0i�v�60O�1��D2�0���x��L^9�0��R��ռ�k�l�F�#H�[���c$'��^��f �* Z^����/�IBR�}����M� ]���ϐ�L�z��n:O����>K~���'(�m�A,�c������W�0�� |������=�Sa%��Bu��B�O1`b-&��'0M�|\�q�-��.�Mpp�;���X[+�!ʜ,���\12���O��>O�]� ;/+O��갽�rXS?��X���w��׃D\�;�?k��<B��$�p(1�ʺ�����*��L����66���Kj"Gx��$O��|@q�:��!T��br	��2)<���Yg6_6���D���K{���3�7�|{���Xr��?*)���YI��j��������2�ĩ�YF������̍S�ü�������;��}�9J�O��|#��`Cd�}���6v�H��Y�\�Q��xNMv�9��ܗ�W/�}�[����[[ �H"�.�*h��x�9y؄��l-ޠW��aC�ƑE��dD뭚;Z<����V��iȓN�;�ˬ���έ��6��.4iĐ�Fl+�:7y*<h��]�H�5�g��V�&���}X�������O}u��
E/���_����[ÝǇH�
ze�ҽ��2��Y��y3�,��v�C�3j2�wN���I�C2,]�hE�y��k��פR�3�.,��-)lh���tQo�P�4~C>�g���!P�	�U)-��N�BnD�u�H[?��dWC˚\@xm���"b�5IF��'o�!����^dJ�~'*(�L
Ә�n>����7z��m��_ih����n�m����%��N�л̝�1B]��e��^�LMmH�R���Ͼ!$9R����/�N��F��$G�����<Ͼ ��yj����!�K�,����[�qT��f�����E+6��0��d
��ex��B�Q�Ţ
�D�U5�ooo�-:��J�W״B(C�|�-������)�(���eU�'T.8�g8z��-���Y�~9SZE_�����Ө	F3=�Ew@��;�y�_�\U��kG��K9tb��Ǘo}���P�}����R���<Ly�Y����\���Q��W��Q�q�C��s@\,��B�9ӂۄEʹ�\�a`G���#�ֻ~�I��s�_�L*�l\�ީ��G(���s!��=����݌���j�.}��ya�P�Q8��hV�a���}�8�m�Q{� Ǆv�2&�S �u����	��斞 qR��I�/������,lmў���Y.�5S[ݹg^�������s�D^��Y�;�l|�ƪ@ �$�u��.d�f��F�H��d����F��L����C���e$@B���:i��z��~���[>d�<�q��H�i���Fs�Ιi)���n/���9fk��邟�Cd.sN��+�;4���X��6���t��^i���D͘����I�����њbA��f��H��lK,L�hjv���(����N�c�C� aX5B۽ď����=�^1B[v����~���~�b����M��LK�*z%{Z$c(��߲��d轖Z� �jX��.I�X0��!_�����,�Z�`*����^\3U5F�a�K~;Nܜ���5|�cn�i��X��m7�	��$�4~���J"S"ިp��y�;��b��e&<�*�1H�G r�p+{4�Y�
O��
��l�*��Ь��֣h�S��	J ��Ŝi��`�T��}����F�@�/����{��X�_3���Xj6�&۲`;0,?>!��7��X� +a߄@t�����%��#�.R��J�tP=ч��2x�[<4,�4�����O�	�
�["�@��V]��n�*^���f+�1����i�����pŷ嘆�4Q��X�T��M�54~���3s���E�-�D��:�1�-դ�F��E� TA��Z}�+8`�D�d��W}�> �X(�/��Y2���^�s�� �3�I,����n�U��l�_u�c.�br��?E�����C���F��n��5�C?��)����P���6O��/��7����\��-��	1���o���g�j���+#���Tb.��f��ge���t>�#ZdF�7j�a���Ӣ��DUp)��L�G�m�\A��F�Y��٤րw��-@h��?T>�P�B��������Ў#���Q��,�&���SB ���kD�(<1�����j90�ݓ�mvN��I�z��]�B݃����/"��S���������AR(O���TJ���^�Nx��.�j|8��}��~tXW�G���l�A;+�P�~B[�I��6��8d�X��A���MV�Eâ�O��W���)s�J��<_��#�� (��?5��fbz��'K=�ى��=L��H��ˡ����ip�u��1�	u� 
 �e8l7�ѕ#��Q��.��`���ovv�w�\��ᇪBL֑y���y)3�q.�&�6����}��OUҬ"; ����o|[���	��b���cԾ��+�"��AQS!�N��4v"��\�J�\��$XK�wͦj�E��+iq�P�Vs$z��{�?���3L˭�dCtRC��_�d:��`p�$V���;(�����3�m��a�$$-hO��}5u�Q{����X]�i�Y��������j��� W�
�8�ڜ3o���*��>����:�i��맖���0�7
ہ�'Uj�Q-(WAf?���D�3l4T�����:G��F�6x�pw��Q���ơ�$ˀOf���kȕ%��ӝ�!
l��6Jc U���F�E�����BD;Xqh�XEk+��;��rv�9�=F\1��1���#�
5\�q�P~�7��/�ik�1�n��Ė}Ϻ��w���2(�8q6bO�e�̸�[�lO��y��ӱ��)>���9{��ʁJr�V������/�dҔ� K6�jW���H%�h7���d�X0���9�T�������9.P2R4l�ۻE6��]Y����M�/.��p�p�Zmv���|�Rdu1i�&�����X�ʹmF�~��h��`R��+��L�H4���S6$�v�Eu>?b2�T#�`U#��gb���Ɠ�.����<�(���~:ٙ�ׯ���%[I+&�^G�J�`Y��s\��Mp�v�ǝԧ��X���po^H(���@b������dl73�j"����6+�Ih��
R��j�Mo�|�)M�c=WH�rGގsQs�_��0�&tb��ȁ��� �(�u���G����_ē�5���RgnO۸ɩ�&#b֔-��5�Çs���^4wOkx�_��<ڋ���U�}nzUM�v3n��{�|��E������y�q��$6�d` �]��l�$���#�r�@�3JO2��P6q�r8V��@�{9��$4m5@��hy�Y�Q�5�_4�?$�ƀ�ŏR�5�n
ڛ������r�#�+Μ�-���U����Ir�7�����D1o�@2���HnjX���2S���	k�D	� sh�$��m�?g/�J��x��S���<(��P// 0R�_��i��im�\��K�/6h�rM�r�����������4�C�xҮ����\,6�$�j���*�(>�VP�Ԭܺ{��k��:�&�q8]¹���W�P[�h�J ]~0"�Cx����a��*��l�C�. s�@���&�g�������}�l�ayӴ,�3Y�,s��ɳ���k��t?Sh@ǣ[�Ͱ'��p�>�Bmgr�z�&���ވiX��W�x�0P.ſe��5�]��`�N:���p���_�]+'r�
��Ί��ŉB0���k�����������٦�aSt��[�������5�*¤��!����'����CPV�_�es��%�G�vɥ���PJ�C�GM�u��7�F��b��]���"HB�$��������R� ��\�"՜���'�����P�t�.I��z��3{"U�9��D�_ɪiy5����,9���[�?M���ma*%v�'��t:��:�Ό���6e�]V�¦с����ttq#י\�y$�t	{���
�\�2��F�p��:��٨����%�B5A�]��C2�<H��R^��2KBd�st�%�9*���ʷ�@������\	5�?�2,e�tj���8� ���=�u@����1���^���c�R�X�وW��t���*��O�=;6�ߞ5!o�&*�v��ΚP��~_sR1���9�F8}��U���K�5]߷��	\�uU3W���#=�PPC��TB��c��m2���r^k���>DOf���<�@iNH&�\��Ff��Fi�Y�@��ټC�,n^4�(� ���p)7wL�L�ݷ���ZC��78��x�}��"���c��Ƚ�c�j�Z���BVH7'r�r��靫�A%U>��?e�� ��2�}��;��Qd_�j��&��E�c�Y�YU�Q�1����T87�:�E�Z��h^�����0�eᶾ'��jUO�tP�P�� C���e��h��=Q���;�=]��>�	�Ye��qF�[�	|���D5 ���]�|G�s:K���|���T�����;��V�-ȥ�^$��0W��2Y�0�h �7s����������
����R�C����4}�#>��j��V鹇ئzp&�'U�&�3�r #}G�Wv
�MNu�3*y8J��Y`ƹ}��u�$;6��lotW+h.ev{�AB�E������9�֤�F�g�mm�;!D_Q�o�Ǌt8�l�q�_6����C��xO��p�FѮ��?��~O����Aʝf��YϹ&�)�Dۡx�uL��E5n��nx$����[���O���#PM1I��yF���~� �k6�*�aq��ä�c�j�H�������IPڣ3Q�y*�ٹ�80UZ���N���@����9�!̵έ���Ү�ӸG�a��CFl������X�����߯��!� ���u�V�a��@�ᚯ���@�'8��:�i�|��8Kf��FE�TLҰ:Y;�+7Jj�U�(�e5��.���泽����Hh6X��ڳ,�Ēg����ˉj��ˆ��]ԓ�T�b�GYdR#(��Eg�F>�MC]��B8[�� �'�n�)ͧD�Lp6�(y(��3��X��g'��h��CW@����z�j�`����@jX�.y�37�zSxZ��O���G�цv�wͮ�0V9��h_�ȐT�>.9�}9R�T0=��Y��3I'�VX�PM��U���� �h�t h�ğ�C�ڞ1z�j�:$��P�r�+��i˳=��)��r
�fs^�6[���v���M<Ƀ~q����d�`{<^%�=�o��������ti�	����y�9-��e�(1�I� d$��$��̽38�bbhqo1�ĳ�@xF%]�6$���\ٳ�����r��BlQ%	��Sc�`��?׋�g��SV��@�;5����j��=�MT6�uI�8����Zs����+k�3Y�	(�޶竰E���F�����bwݳ�����?6��e@ Ff�"�<ٶ&��`q�)ޢܲ�Z�c\�Q���^�$iωW��ÈQއdh	H>������&����O)1]�������
P���r���r��`r�y�ӥ�dm��}�F-}im�2�-���dL�_�M����-�"r�G�I�,����)��0F
%���A���Nʪ���z���m���kR�#���>�*�Ac��e�vjם��=hٙ*ٴ��J��PL*�5<� tՃ`�]\ȑ."��h̓�˔�*tL��(hA8�=|=��no2*���#n�&�ڂW0-��'eI�iB� d�~�� ^�z�!Y�C�y�e]��sُ<=��`}�U��w1���OrF��&l2��-�.������㞽��}ݩ�S�,[I��d��-�'v��:"A_��l> ;I�7\~���L�(��.��.>�ī�J?�w��g[^��-�"�j�\�,���M�CSr�k�V��
��M;��U�t��)3�Ҕ����L��?	CaE��?~���B\趉��\�8`���|�?��AOת�Y`�R��a�K5_]��7W�R���M�$Kt��t=����_ �z��܁×��q�{E_�1#��0����D�u�֦ �O�1�ݺ(:6R_�a8���:��6+ua�<�� ��U��UNƞK���fM��;!�^^��d��qD�A��<���ʖ���ɜ0d�ʐ����64;FD�<
h��,�1_�b�iO*�(��:�h�*}��?��k�����	�t㑹_�{:�%!�/����[_d��'Y�m�5|��\(��u����L 
A>�p J���ն��)�T�]j��PB�\�v�J��� ����?�t�<�4|���S�ք(��(��6_�^���I�XG�KR�Q�ma��%c�!iM2��F�yr"�+ ӷ�N�)}����׉� G��d��uˬ<Jl��u�g6r�AX�r��}�����0�C5�*n� ����Z/8G���?f��P�x`�[ح^?��@؅�=�6��l��Q#Z?Hr��ӂl�&�/�r�2c���[��aB�َ��>�2w�D
�e��l��6�:����K#�M�om�\��Da���T88)�ރ��w�3GQD������^<C~�MN��̻TzK�R��������t���.]%�'��\�����P�}���{l��K .�O���2�F��iG�}Y�S�y-��c'�f�(g�!97��@����A�xE`)�O���E>����_	G�9\gy8��JE�?���8�:x���}W��6�w,�{�cv��H��΀�PCﻣ���[�]11㏱���.�O��!�yS��r/:����]�8�S����<@�'��qo����,"�B��o� W�h��E(�$@���?�Ì8i���S�Ξ�2o�LӾL]�y��Q�.d�����t��{���l�&� ��M~2��=y��2��?�f9f�.� �1��Td���>�d�X$�۬�7���d�M�>���n�+4�>�	�E8yO��� �c�tK�8`���'ډZ�gsK��/�c���8���^����+����?���m
.�1�����Dl~u���a�����蔰�� '��ܛ\���H�2� ?%(	�L3��f����^��yOy��6�V�Ȟn���~9�?���)��#�����bT�+���~2ٓ���[dP��1����{������>��&����_ŮDr%�����_}��<�A*mP
�%�Np?&<���h��vK`��ص}��q`@iN��u�Hb�D`6!� }8M$J�C|}|xŻ��g�7�r�6Т ĭa�m�K���TS�%t�u4��W�L�]�=�J�$��uz�Ǩ�ļ�@�n�k��H$�a���ra���7}-���!?-v�\k�����0$xt{ n��=C��\��K)U�D�����^ӏ���[��5��+������;��AS�iq���dRL���L~c�<��{�x:�C��X�I�kɟ��аi6�jݕ'�`E�]֜b,��R�����k��a�]�-U��
�UIO�d3��Y_>]l�$��� ؀!�ؐ��joisF8>А,&�w���<�����)!g_�Ĉ���E�*9a�KlJD���j�^���.CniK����w�hb�Ô��]���&SCg]b���4�����uR��ʟ��qvQ�7p��ֆ<AӉ��݂F��"��/0i��A{���R���2j7uԍ��ܩ�q�G.a�������;���a�:����09��L"�u� ��e���e�
S8dێd;��a�)�]��?�#ީ��?*����ɮ�m<�-PT�>}��6���V���O�'����kL6�c�y���'�+�1��';���w�)�r�Y��ɲc�8��m�#�v$�ɘQw�Ϣ=#uB�Wp�m}�e�]�ȷ.�mH�/"��V^\�{ MДJO�H�S)�d�D�4������w)#n��گS$��*�+��MU`�ƆdO��9�p/+v��G��Cj����3Mr
��{�}٭���Z�� lyƧKЈ�wP��.�N�&����r���e>��&�q�}��=0h�ԉE)�����b�.@�hb�7����j)��℞"C�8'�����J��%
 ���ZsI�qR�����
!�����u����~	��7x�yp
���v-��սisc��6���ĒQ�ʛ\��'s3�����91�|�N�{m��(~g��Mn��@?j��H�ǡ'��2O\R�O���c
�
�k��Fʫ���P�8X^F���k��-
]� �����ɋd�����l�j�;��XIp�c �^X�S1����<�`�e���""��6��u��̞��"4�L��ʏ��
��P��b$EO� H��h��M��<��J��[|'��Ln�����d�v��Ȍ�<ޤ��V'b���,����;c�ew�r����6�Z��8�kYƨx��$�1��ՊR�ڙ�w��������|%N��N
�;�m����=���]%T����S�a5|���X���3K�Ͽ������.�8IË�+,aH��� ��l�i?h�����+<�~�A��>��R��7�z�R'|U4}���O�8����f%����/<�q�Xa=�^�J2� �γf�Y���K����쫶�1t��e.'
e���)x������s�����c.�k��C����nn�*^3=���Xk�S�,'��֏h^�ܟD'%І�p��5&���':I=Q	�T̓ŀ1��z��;�8M�oX�{S�ef}ɔG�%�A+֠#q����#EU��t2H֒QPU��;�;*K�e�G�[��o1� �p�?@�0��pg�T�\�TĠ�i,�qP�/��?}ȵ��-�&�֡T��ʭ\k[��:	J�/�H��!+���\>�[����� >� �0vMOY�R☏�[\�j�>&O�y��>�5r3-��Y@W�(� �P|u���>����I��0�1�����b1׷�;M4�Z�\������pq�o��v��I�� ��;�/_�����iV�C�7(���_�h�Y�s�f9*k��t�n��է6�����]6�̟�5a�z�=�}��5��lC��E�O==����_���	����&fahi�e���
���>��a�����r���}ŻK0s,L�0$�ܾ�-�6�D�9����l��+������Z'�X��<!H�;&�����*�##���I��� �����*�Hf^�f���1��,P���A�a��=�	��2���j:���އ��D]C����3%S��Q2��[" ��8{ ��-1;�O���#�݀�a&�~�P<��6]��D��;V[�4%Na>UZТg�ӻta�,���9YR��D=+F9��E�1rɧ6��G,��Mb6�\�{;*n�.ӝ�-4ĺ5��`;O�R�t���*����eh-�X�2r�i(����ޱ��GRnM#O�Ni^���d�66JG�����X~G1��P��C��s���3~A.H�Y~IXi@AFyeP@ȩ�%��xW�Gy(̤�	��Y:{��ݍ����had��3��#���T����=Ic�~�r��?�
�e�:�i=�^LFM��ud�y얯��������}�\���#�:KSK��.c��5C��Y|�
]���¿_��t=`AÿT�Q8"~���"����{E��ej�9H�}!�"����I$�I��V�8�Q
,X�@�-�xg[�M GL��0����V��*(�_d���4v0Մ�`�z�:-]kϦز�!|�#�^Zv�D�FpA�	���m=�.1s��f��1���`��ê��r���v\��wp��,�����(�zZ�����Ƹ�J��=~�b���ɆV�� 0����+`�G3���Ng�1�qx;�=�B}:�jn�v�-m�Q:��zY�"�a��Jݝ��/�_�,|�!J�j��uI���Ri;7Ė�.�"B�|��3�!�� �Q~eZ���������w��*g�\���x�V1�Z�~������ѮG�@	�m{i KqS��¦.�q�X���������^ҁ��)��?�����17_Ǳn��B^d��)�7Lϖq��-Ie�+�I»w��5�1U�W�e�_,��\�?����� \���~~4\*t��5�9M�d�����m�_����E�q���O\k�D��6�c�����K��	��Gq��eVq�cIcM�T�2����%�h&���%^}���&Bǈ�]6�6*�q�)���Т{}R�1�cV�6���[�K�p`."zu�M�`ԟ��9�ʬ��A%#"M.�3��Yt�!��:�ԧ�F�\A1��9�5.<��=&�?��nr}k��2�x�gVZ�.��#������\��.����%��A
Ϊ��>�O�Pm C�a�s�Iv����O-ә^�6��Z^�|B�.��B�95tp3� H�ڬ����N�(�Z�t���x5 ��v�	)��t�3���X�0��.7�&���� ��~��u5�%-|�f�ֆ)��4_�\�G�D����PS�b���d��"і�'����*#O���0�����ᕀ79Mû�l�bj���%%����M���q>���랜���[����ҵ�4$�~"�I��i��9a��}��X9�	��5^t�'
}��V�bV��h�)W�Ϣ�o�!K�E�;��Q���P�F�����ޅ�s�P���jw�Z�?\}3$X`$�.��������^-��|�J~��kM�o ���Rpݶ &�S!�>��C�2{d���\�ܑ����� M����A~���U�y������|O�����Z�K��M��8�͡�~F��hh�Yp�Ǽf���W³��������H� �w�`�_�nN2f#!��Uo���#�<�2����a���)��!��Ă�H#�Ǉ�h�lmwD��x?~�ӓ=NO��jf'7�~�YA�#��J��ԫā�]�fY�Ħxg�H�K�`�O�/~t��,���uWԩ�8�/����І�$tkf�mn���)��H+<j�ه����>���L�qi��Db]%px����z��,��B#S�HY��d!��T�|�u����R��4�6�HEq��R�%����&�A Oߘ�qW���hJ7���{�A�����UԴW졁p`��
��F
���j�d��,d�����E�^>�Ѻ��X:n
�dp*w]*k�a�鮵�>oV͂��~���_�gU�|^ܯl	#�W_��E+y"#�\�oGg�[�L-�t�䩳���o%�Z?M8@�HӺ2�d��4��W�v�aP��3J֟ ]��s�Ќ��`8D��I,-��<$����!X�N���8��A|�rG�P8H�p0Fc���|�2):�����)�r}AӘ2��{)��[a:��>R't^0}�|�k��T�a���%;M�]S�G2��z�|�p}{rS6���l<Jo<�;��;�KL��+��,	j^+�}� �oL��SӹM%T@�	뤏E�@�e=��^"�\q!T�!�b�4�+P��%�6��#�����מ/�^_+�F���a����h0��J�(݁��݂{F�\��r���1(#�����7_�O��{B��
3Ć�z���<�l�l@H2��w���1{�k��c��[J��V]�v�
r`�t�/%aA�Z�1���ݨMD�Ns0���сðhE����V�Y����;4��	��7���⫮T�O��.7Ğ�D���4{
�w�ti%��*����:�u�Z�3�e���}����\A�To�N����<��)��1Z��ƒ��bZ��Pb;�e���euBw����Bų�Pkӎ���Z�13S�!���o���q������|��l69\剞�-E���s�ϧ�(�8�&y��b�#d��oA���Ns�8��Jإ3Y�>�80j��A�y�*��U�6��
�h���C�������\E�GI�f�b�:�l�g�����ho��{>p����1j�7���-H-�¢��O�"��ui��Ț;��<�\i�䙥�=O�I���5�;[���a�-�����m�VG8�g�1 ���	����/��M��A�-�6O�,�����܇�]�i ��Y�@)&���a�)�J���^�uo�+�C��d����h�0�J��Qh��!.�b԰�A@ TjE�^�2����� r�$��,�"�}G�G3��l�E�3����v�]�Y-�{=o߿��\��/le�?�2g}+�N�=���Z}��
�%��Ȕ��613�]a=A�|�KY�� ���!Q�`re-Uy-\%�rY��TaXj��^���	Y����#̧^*\e��9K��h��?���!�eԮ����X�p�*$��Hwg�Uj����T=5�{NM����˯�Z"����S̐���74��k���$��Wq�&h_#ٹ�=��[���/芟$*�8\��a!����|犎g���N{�`i�l�܄]�
�m��T�
w��9�%8"�'����sU��R퐣�TC�q�G�ea����ܼ�LŸ8�������ɍ�JgO4=p���j�&�S�jx�$!!kO�K7:�%�ߺ�D^���Uk�U�upN�F׶_%�h��S(�"�#4�
>Q��	MJ[��F:8+v�#�$��X��o�+�)
��2�R���*Oʨ��؍���R-��]29K�g�÷�G�	O����&�
��]��A�ߩ��3��C��kF��Zm;j�	=�F�o/�;w����ԍ�ߒ_"S�s�A?Z5p#����� ̄�;;�C�˺%pLmcw'ɛ2٨��Ls�!���6��R��ƪ����f�/�Y��c�R �s���T[��1��-2�<�2��K�="/S� <�m��ܬ�8.°�B��O?;�A�cQ�U�n�R=ʭe��,�f�R���=rz�9�����b~�h��� �1�	P	0��Ӧ��s|�������dJ��O���(���f�x��\���pzD��W�4������S���6�:�/�G>N� ϓ��(?$}�G��Z���5@���ʕA[��30���h��k^O>�6����pzX���%@�����rT���u�؆i��t�;ሒoa�� ��/�%��6r�gW$$m��1W�r��cx$U�B%Hg���|9�p��wO�A�Pmi�4�)�Ul�,��c ���o�7����4�И����3��`�|����W�@~��nE��.�o1AJ�~��x7͘��:rF'�Y�-�Z�܎����N���x�/�y�K�| <!_HMFI�O�cE�������g��v|�6�_���b���p�X.�`��� �1	w�i@�<1�55��ckWgX� ��,�;�F�V,�⣯���Sԟ'����e���y`>�dgoۆ�>�~NdLb K��m
M�Z��w��u�&��Ƞ;�-�x_X�R��JQ�q��)ς�u�Cg��䊯��<��es��p�>|���#��'2m�_�9�#1��K��ẈG�����M�� !���]��L �%9�=���餙W�~�r������}pɢQ�hf���)���A>��ψ���98��b�4�$`�I�t����F��c��ˌ�(hH�/Br=D�[G��B�����p~o�Y�W����{�P	��@7�����ޝ^.7T�!�N&�dF���x��\������\��"�&Wh�	&f����#�W!�؜��R�l{LY�O��)���T�q/��V��<My�4g����3{���W%V(�s�ʅ6N��4֞D �J��9���#���X���L��Mδ�{��s�Z{ĩ�?�7i)�%+�@�*��m�MX�{؈A#c�o����@�M�RYMw� �>v�Ű�x�Ѕ`�F�mc���mZ텀�t��C+Y6�7��<��rCs23�Ę��J�w($x{�| �)�i�0�F$��CV����;ޫ��bo^^�;��)�br�J�Y&d�tY�l��i�I�����֯~�Ù�Ӳ����l �X%^Y�����q��(�c��M;�:���/�-��W�1mW{�N$�Fa�FH�������R����W���6Go
y�������n��R�i#��%¨���}	��F�z��g�2T��x��^��+��Lf�w�`$�۬,�'K1(��i���m)!�nA5�z��~e���Kӭ�ZVFwQʰ#�d��O��D�y��w4��za��&��4W��2�P)�C,�#���Ob-��wp�^���Tp�U���N쯅��fF�/�3"��O�s N��! w�F�x7�#�z�ُR��"��	PyH��2��E;�����'�]�`0ǊJ$�=a&�^'��d���3��v}jh~�&���q2A����7t�\*{ g�]�hA��slb�\�f�[����6�EL�y7����'�_]o�\3uKm��ݎ((`�S���h�r�m�Ҝ��7>	�	�; aC
�:ά��1@ۦnA�kbg~k���Ճ}ԭר�{[�g�R^��h�n!򾳓zO�T�������U�/-���W��v��O�$h\3d�Vr?�ޒ;'�O���H��ܗl��}�)}��&�g��XSU�ܳ�̹��e��,�p��<Ǵ|T�"�$�CG�p?~���Z�UPa�=�dPbw��$�T<���)��IHXŇ\�����$P��^��QE�5�d����ˀX�i{�	����V���.�wz�, �'��@J�� ��疖�/o�����iF��<ڼCK�o�J��T7�g��|��A;Xf(U^�+���(R�"�:p�"����R���ůrP`<VA������
��?c�6�ϒ��s5vc"B���R^���������m��^�b]Ц��`�'�pF�5�:m�[�~M�X�2?2�����2ZvS�m<�)�j�5Íƣ��%��{�ŌY���5
7���m�	��}��d��,�i4̊W�AZ*@w���$�J�h�L_���B*\l]�O4�	�iNI�R�V*���9�������,��(�q4]�o���n	��I.>.�C��#m�܋���(�o�!Wݠ3e#A4�n�	p`���؝%d5�xp��_`n�&�U.2��n�l�.�?�r?��
V;�����7�b��J�����fC�t��Oh�x�qW�˂eVqf�'���6͔���P�Ƭ�Ur3_�acr�g���+�6�D����bw�˭x�-R����7�ڽ����E͉�#cM&�g����<�v��φ��݂�����,�� a��\�l����H�~������h8NEӉ�2�0d˗k	��5x.�z�aE)�`�;�3%&�&�=JH��:�:\�j�&^��
s�����V�?[�+��$w	�fMO�$�],��# ��`�D�/����$��6�����x�XLd>i��A�˾�m��Uo��Nl>+aKH���@i[��4���$����T�uU�˜���m+[p���e��1O�9A
yko
ؿ�D�(f,J�\Y�����#~�e��b�;��\�>�B�� `;N�g]��t�"+E�S�*�;E
񷚸�N1"�;��7�&�q�ojcťO�ٽ1E�5;��~#����Lq#�� �|�~� ���]~�q$�o�]��Ā�zڧC�9�K�:��^�T��V��V6oD%�$u���*��9�C��Moc��-�B���ɏ���y(g#��")/����0��?ŵ�b���?�K��OP}3�`�揫�53X�KZ4�t"*�mQ�G�K7�=���:�X��n10��0�?�/0)��.���d��;C`U�
i4OSl�[K�wZ�7/)��p��P���Q��<!FèJ}�7��R�J�|�qO� _��p�l�T}�G�9s��_�Ѻn�������U�1���H�c�v�Z�B�閴t¶���6�ȱ9����f�.3'��`�C��">rT\�O�?f�d�b\$PT�̳�Aɛ�gu��� lqsGJ�2խ��B��G6઺���gN&^�76�zk<#/�RJ;���j��8F�`�Q6�+�o2N��E}�ע�X�����DU������Wg�c�!ϯ����qY�ý��R��&�<띐_^�m�j�nBX��z?�zq����d�o.I���'���D�*nW���I��7�,�]W'�V�x��QN��R��&��X���k�k����鏔=p�3Hj�¾��5��8H9:9ʠ�JT3���1�o��D��ǰ%��\ۓ�K,B���O w�����,fA�7�j�$M������Ļ� �?�E-L�ϒ�ɚ"1){)s��n/��#���ot��oN�R���u͠���H�V��|(���R��x3�K>=��,��J���xT�4�7���b��n2s������7�SAla�4I��3�%���;L��Q�M�[Z�^�E�[���o�2�5�Q�DVk�=n�Y�łcQμT������פ�G%����iq�p��:0 "�b��eZ\.��͌e��L���B$E嵚@�gQҘ��3��uf��0�zïw��~�p��+l�(��3�&,�7
�op�-�_�� \�X�����<�S����l����<�Dϯ��@l�>�h:��Y��?ȱr��JG4�(h%��e�-tv�p��A�9�\}d2s�}������2���A}S
d&&�tP���P:o�vGj���D���ͤd�:<�Q_o`2���$��E�s�y��tHE�B�u��r�1�a�� ��B��R�IŨ0��x�ӱ��MZ���]}��1
�	��Dޣ�bկL�)��S��б{����T��8rCt%j-|���sw�����s��TfM���$,���b�q'��8>ZѴ�6	�,#������n �虁���'�v:,=xk8:��l3o!���nx�Vjr���\�Wl�c�^�Iԥe�����Eh�v��[��h�T�Q�0袕Re��E�}-��U����ty���_�,�k��Y=�"|�6"���Z#��l�K�lA6)T�V��ڢ��]�=r��:��o	s��4�9ɉ���=�4�0��ks�����#뢯��.z�%��q�w�4�MG�?�B��Xk�3��>^�c�>nv��w�(���,�`��]��wrx��j�_��I�$�����5�A��χ��z{��Ĳ�J�ۀ�b�ҋ�-��ӤZ?!����&H���YS�g��`��|s�Q�����l���\ȇ�m����~�|��:�K�m�3�\�}��}|�g�t��_�v��o�� j�Ũ��(��:NT�esp@f���\Q��׳����㧜
���ZԂ7V!��Ҟ�� �.�#�&��O^�!�dz<p
�ӓҳԨ��AQ�$.~i����΃	��g�iQRwu61��ߍ�$(@%��\���0�ٕCg�-��b㡚�E��C�eM7�َ�Ĭ��7���̓�q�Ե�\�p�7޻ڢ�?KT�k���7a
b~�Rr2Tͺ�q�rP	Y��_S��	��V�b����)�Z�R��S~����v���qQX�r��L����@��7)������nW�^X��Z�:�<Я;q�UZ�A�N��&�F�"��Ny~�!=���,+��L�u���-���1�k�gw�$s}#����BTn�ҷ� u�6�]d��ā�
�?D3��F�[��A�φ�	�Y�z���Q� ��z�*�z5j��)U�Hf�z�O�(�ľ	6�'d6ܸ� ���7�%4U)Èƈ�%z��K�\�BA�_��n�x�^��7O6�S��-Z��p��?����Ys��a��$����z�Q�mO���?����1�Hʅ����p��y�+�@*�B�<l�0��=�bJ����w���;GF�����k�R��-�����Y ��i7'��yV���E�7=*�8���I�&LHt�e���o�r}(r��Xnx�gi3�fT�����@�������BN6���g I�_�@<���sq��?<�����Ƙ�V{B���PS+~�Oe&�8#��u7 ܇�O����nJغ�C��LD�����%�ۿ��"޺�/�ko!f�<6�����i\o^l�["�g������%���;�_  ��b��X��/���Y����t�8�˗X������=��S/�d=q��⡁D�������/�>l0����^2~'9'I�Z�Qq^���Dq�K�Ls$(���7oL�4=g���QG�8�U	�aɔT���)3g���+!��~c������}[v�Ek��1f�8���6���z��ݦ�w��28
���"�s䣈x]�NX1�p���gX�A�������͆ �dx n�ŷ7MW_ހ�M��,��eƹԩ��Ҟ� �ch��¡��"�ڂ��1�����n�� �J�w��v:@�C(V(?a742�x��/�I}$�]�B>��
����w��a��+t���d�DJ/����[+i��g��Znm�EC�p/%��>P�Lޞs�� �䛇�=�VR�S%���{��O���ũH��kY��5<�1�:۴�W�"����eP$W�i�b�� ٯ���(Q18�qI{������.SR���ВD�a�O�Ř�^3@a!ed���D	��)ъ`���G4�4�����*x�H��<���T�XvOkٹɳ�H��7{���4��ߍU5t���cwj����B㧤Q*��&��vD�r��Q����ͣ�1�~ĩ:���l4�n�ζ��8�b�fZ �_o�������P�e��{E!z5�4�:45�� ��+{��(K+ �!�h���ϖ�6��sM�	��8(ܯ@�X �8��YN�޼"V�d�n�Q���n��\q�	������ʍÉ�NB`�e�*�,�us�a�u:KZI�+X��NO/�p��z,��M��G!��ɼF��a�a�anMDk�@����:�;�c��>�ݩ6��N��3x��m�Pr�A��_ �ä�A�>��npվ��<%��J�;5�$�":xo��!8�@�Pc���~�L���6��8�̂)�4&�N�\�=�Ux|)��)@<���/S�R8S�$@��y�QEc��_M���ⴒ	ɝ�_��H�f��Qɖ�	揞�Q��.K,nFw�1^��4�-X��M���dq�>>U�����L�h5A�0���w��
��,��O�B��R�x�7�����ʟb�GrCe/�fA[w��G�B��>G��9[6�:,"��i���sH���>�����Q׍���-Ɨ�;L�2�:��@V:�+��A�i�C<1�4��2_���TK��h8����Q'��_`Gz��`?
��R������l�@�	L�=6[)N��}�X�p�5�#�\��H�te#d�6�Λ�x:Ws��Al7f�|9�
6�3�4��ĝ�p�f���x���!��<�/�[���������>:�4�5n�kD�7��j��q���]6� i} '�S]f�豔2��8�>�Ǚ��o�)o���t�f9����6�iu-C���!v�=�C�x��O��e~	UִT���3�#�\�%'_��'��a*�nd�w��~��2I7�}����N~L�R�0zt���1t`�ueR�E���A���C�8"�o.��N�}����9G�n�ZA���O(�1��i�+5��q%O�(BN����@�r�s��z��hʎ�o��$zU�h`�nؤ෬t;���%����號�oƾŮ�ԜW?ܖ���m1Բ}#�]RZ��'�9�=`dO�D��%�%��"�"PZ����,ۆ˽೴����"T�`N��Y�������6Ro���G�9�2rWˈ�8G؅�$��,f.8��4�s��U�B�X���(�, �^���;�$|�
�2�q�f�]D��3"Tҋ�(�Ϙ}�(�w�1�Ic���xH��ՠh�)��'�gͧϤ3tF5�/Ƈ5-wa&|L����~�}�����$*���yc'��l���>Kk?�`��� $����z�0D���W���)�2����H!�Hld1�?����X�CEJ�GE������,�G�ҡL+8 `�K�j�F�cʣ!��e6suPS%���i2���i|ׁ�N�G`砱�0���k�%�ȋ怞`�������sS�E�Q���@���a�Cna	����I;�.�Cp
��^nԥ
AQz�ִj�������+~	֔����X~��GĹhr%�춣���p�v��N�&U���%/��zVp=�6�k.�"bsYrF��Q��������B� ��I0h��Y��e��`H��/m [�/��gYT���i��N{��O5>�\t`�7��zo�����@D������>�$<¿;N�qW�:VE�'��Oc��UD����0���d�n�,. ���Ǚe.���2��u�!@s1����Yc�+Ʊ���{�uV-���^�c�c0*����N��n^�%�9��fZ��@9N�1��Y��܃����Ӏ+ю���\H�����<�5N �o�����qX�p S�O*�R�3�o��ɐ�Ũ��瀽�4d��0�5�)q��9R4xJL���3y�Sڝ0��aғ���B��S��Ԩ���Y>������ꘛ����	ۓ��\}�L����YN<���z8ڦ!K�4�8]?K+��1u)�����"�D1��~0C=z��XM��-6��m������{��+C<��m��7/�l�q��`D-��[ѷ W"L�)\Ȃϙ�H>�')W#/˥��;�X��y-Չ΅�?���)����H	��E6uj(�}v�R%�lt��e+���`�6�|��a��k��g�+	����G�o��V?==�8���b��Ǥ~�*)6�����B�!:�����i,h;��G��й]Bs-���|�K��#m�B�Ǹ�i����X��*����r��,Kō׶�B�Ѕ� ��]OZDEx��7��27Xq�e�\M�ن��Y��8�T��Q���̼��M�BO��X< 5�p?��p���')���
�J[캜�����\�p|y��=LG%�GrƱ�Q����9��[&<�V%Jfx��Ԭ���~����g�z"��y-?���Cuf��!�� P����|�|F*���%g=�q������u�� s��܊�Ҏ�u�7�D!���z|�`s�D1��d�ǝ�N*Q/�N
�C�vv#���@�Rh����H&`��nػWF6�)���;�}Ӄ�b�7���/��4�4K�^�!酻L�t�A�4g�6�p�y��c�����y-���BkN�L��1���V��~Rѳ>c����W�:`�����8gI'��  kI������es�vY�������F��d���+*��з�uZ��,q��Z[�?����4d9F4��#Lr�r���4ͅ���ݕ���,Ԯ�[uEh� �L}LK��bxDK���q����q���wi�0�q"W� ȏ��D�{�o�W&�G�ExcQ����|���������s�H�ڄ|����<�Mg�~ �����A�����4}Q������X��u��k���:��He�l�jA]ʸض ��C
�����1�r1�ٽLp����#�8��C�`EI���' B�k�p�����ڝa5 1h�@>3��͓눅ܷ4������q�/�+�!�p���ojE�fv~�J��`�Nc}�"�����[��;��Шُ;�_���r��M���&r)�x�:	���o�(,�h�!��?���Ǹ��V-e`h#�|��p~��L�	�O]�WW���W�1�ы�+�XA}�N(��!�f����!��=�K�6|0��{R��V���_��������:h���kM���k"�h���y�������:־�(޸h���C����k�>�k�䫉��=ٰ.�:�Ȏ���@/oyg�/q��~�N9@֓�#w"X_�%�^�}�H��1|���<�6L��P�h�4�2�q$)�����ɵ𾦛k�1�����W�J%�^!����6�e�t���C�0��m���NŘ�nO��\̰R���@[U��r�G]?x�8�����J2�dN|�T�*}�!Qa��Z���9M~A�����Ƨ/��xB�ӞZ!ϣ�;K��;:�����Zz�º4t�
(�V��MB�ԅ�v���k��p<&��qF���AZ���\���c������:�B9�ʋ\�ǦZ �~8�;���~�rvdw'{֤��N��/��^�����?2�{Z���z�:�\�*�~;���.HB�D����,�۲�������|ʎ�:��X��P��&�m���t��Db��*���E6�]n��hn>�Z}{�z��\j;��fE�+�����ܩ���b�nˏ\�V~nv�[t���)B��G�$B��8��-?�R
��j��	�_~�6%��6�o�Ą2���/C��f��
����=a��f#��L7%�]d�j� l�Ι�``8��
6[����R�c����<��o���Pz���K>��~�x ������^��W�[�r-m� ��q�c������E+ȡw���_�HM ��b(<Q9��`c�����Ȃ�~鳟_| #�-�&����u�R;��2�KK��~���J��b+P�)�(��e�W�dq`g�e� �O���[y���p��7D������U���ҝ�QY�AĔS�dKa4'wwU�e	e�߂�0���A�3o����O]�P<��%ԣ�XM�E'��b�\�ǈ����8 �l���S�����ƹ{��],�3���+��ɛ�����v�{g�.�ˋJ�� )�J7���=Q+!�፾&@��v��:�Y-�d���xS#��>>�rm��5�9��#m�):a#�Ԗ9.�<��t^�8W&���8���Vd�ג����W��ur��K2�_�9̳4@w�*�7� �q���k�}��bm�3$��Wc��M]7sA=%>f���.�P�9�/����CZ-���v�V�N՘��o�Ҍ�3jX���N�>��Xs�:sHb��� F��8?��-��j6����-��eb�s+�L�gu^���ySl�a�eH3}4N���0q��ԫg�X o)��Z�u\9��,;~��G��V��J�
��v(�����O��3%m�p��ҵ3<�LA�{a�㦙!�K��u�e0evQ���Yh&�	�c�`�kMŅ]ߧ�틥�n�k�c[�#���*�k	&��Ȉ�ѯ����}��4��� o��\m���D�\��|�����΃�ו/b�3�j;4W�b8��nZ�)��]�od
�L
�PUH#q^��87����)��ák���̬Rذ��W~]��},�o^�N�DU7�����Ռ~�@�<�����Nj0���;N@��b����mDc�$�F�8�1�\2�Ƴ��bCU��8����A��y���;�����%W��!�p�DbY��Q�_���Y��k�[=U��+�Z���i,��[J��+P:$ͬ'�M�3_�Ji�\9eXD!Y�R��v�vT���(3w�ɗ,}`�c��]J��61�1O!Q�}����=����a���=)&��)���d�J�հ����=�z!�Ap��g,Ө5���"A�fQ�iA���麍F����wM�Z������+��\c˲��"aGz*"ኳm�5�j/��u����[���6�
�v<����Cʂ�'w��~v1��nE��o̖L3>��|���������+�����Ϊa�x���rp\Z���Z��4]ұ��k��3�qY�=#���h��ǯY7}�L@��T
��NDU��b�����@�����nZh��5|56 � �T'|<�)���#� ���W_��:gy ~y!�MN��SO��%h�������V]��K���d�� �<�ָ��9K�g�VU6��<�`��}I�㫙��:@>'J�ʨ���^E@��r�b�	kÐ�XbY恽G@�H-e�ׂ�#��%��1�:kn��-~;��`�o��O���=u���@dr��'�� 󸚻+��
u���<���%��S�j<�Ǟdð@�n�j<R��k^
�!.��qi��dȼ0���N�M��55l8�~2�4��ȺW('�0 �*ct��)�*��t���b����)�ڑ�&^?"oB��&����K����El&�� �(�վ�R_Q�N���Gl �k�>�3rm�nͮG_2	�B�' �	"N��������A�_��Ts���P�̡2oȇm���E.�L\|,ǜ}�lh�W��@��uZ �R��^�� �\�.|��a�
�q2��+&��lh�$.\`�?$l� 6�� O����B=�s�[�Bt��e�F�v8�BC��k�p����5���o
��}M$���C��(�_hTn�:�l�?_�a�z�h�����3R-��1.��h�9u� �� ���u�`.eϸv��1|��f� ӯ/�I�
��c|�����($���:ſ�	�������w�OQ|nN#{f_�>�&3)i��W��9��]Q%y{�L͟���N�^�U)ؐ�l�u��j�$p�|Kޒ�N�hc���2ɨK"�]��~�[�x)��9�X�����]���v�1꧔z�`����A$0���y�=�Z�Y/��q��_|���`pフ:W���o��`�y��=hY��YV�B����:!�՚.#��GWхll���d����q�v�@�����9�D &�����Gl�N�����'ѷ�9��=�Ƨt����� J�LB��)ʳ3j���vU�����R�7��GsBR
y٢���Q:��U�I�Z��Bk�<�{���g�o�)\��zh*��ƚ�'��_�/H�b����ǴDF�kt��"2u"�
����i&O�k���o"����6W�](ɿ���,�Q�ql�<��U3G��}bp���su�Q�DL`�������܂J}P��>q�d~�[�W��Q S{'.�^�]i���QǏ�0Q�t�xV�'�5�7jӆ���Y�7j�G��h�@T{��\��3���R�V��ȷ��5ǳ2/�S����&�t��������y�*�ϛ��!�n$�<R�tń2N���S�IL��X\��CƦjKf���;��F��C�\@�I�}_��������I3�F�w72mX3��Q$���m�����2Ƒ�Lf���F�x�]WUq4w{~8��@{/و��z���v�o�����?�$ِ�_�)�G��_J�iSG )��ї�7 ���L�k"��7��6k.pq����M`A�E��R�8�(�r��(W�A�7��H�뵅��C�|&�!�Γ��}�c �>T����d��z��?�M�l��'͐�9#Wʩ�{���Bg�zj�g� �Qc�)����r�K�|�����&:	5�u����J?�����Ni�gʌ�d���ɡ�=�BH_����?���+!�P�k�0<Fh������5�t���.��
�_&{�������k|/�bL|��4�M��z���RZ�KC�, q"��0�Ki����ހ�򥻒��.��wV[X�����)R��S���h�����/���s��#&�լ�dgH'�O�vv<M,��ݵ`l"C�v1�i.��=����	���P�v�H�db�g�l�����tŋP�.n�t��J����� )��e��ޡ������ Yɠ����E��bs>��=��Z��t��IqsE��I���s�����l�`�K�˕��]r���󁑺3 ������g�X��賑���e��&�7�qW����5�Ң�������E>�(X o��EIW�5���`�tte-W�!�2��a�$��}s O��0��Ԏ����+{o:]e�`$NEr�//�ʡ���<��U]5l'�뛹Vrٿ7����+͂���,�H�<�:˱����q7W�V��#9�,�4"����q�]�+i��Z�0 ��#��8V<z0R�Nc��i���&D5�KE��T�fV��0ѿ�)�##++ǠY�i�p����_g���M"�!�ۢ�����o�-3_�|m�n���L-j?XuP�Qxz:�c ��N��(A��]�S��ta��.�[�n��lP�����2ӻ����i�Ƀ��lrE���ta����/t��W�J`��\�jбF�$
?�ű��o�M���T�q��7�n^���gCB���#���2���!�XK�OC�t+Y�~E�5z�)�Џ�#ʤ�E�"���2eb�ϣo�A��[M �''�{Ș9��� 5ҊJ������V��D��-E;jɃ��%;�n�d�>t�_V�eX;�B׀}�%M����T�z��Md'��fy���z;��^�ܳ&l.�!�a����o� v߳Ib��>�x�+-
�����U��ȸ�����y�'Nc�}u`�w�\�
^*Ӆ����k�O� �$n�!8�;jLB��Z�#|f׺SP��S�P�y|I%���묥Q�Os����56nx��R�}��j���}Nx_��K�G�RZƶ����h�^�F�1�{��ǀ�8�[���<_�����
N�Z=h��?0E��q"��S�K�%Ub�l�5�a�k���$��a ���2��e���:�B�G���^�QG�wLQŠO�f����r[�G9�����*C�i�X%!�A�n�~No3�D̔�6�f/(�?T���M�ڜs,t �ܽ�k���s��aʢe���Y5!q���7�}vu8B��_:x��nq�y��`��)yl�>G�:}m0h��y�_[!��giS<����{�گ#���YG�&	y�&���̃�.�]�|��<A���0�@&��q��b�#��N�/�Wh%~���dXE�;�|�:�;�܄�EK�{�#�I�P���ȗ�0�b5�W�j��m�gI�K�uy�F-��ql��l����/D�°O,2+�5mC��Ě�ܛ`>5�[��N;{H�������z�+Jχ0e bA��;F�� ��^g��"@K �_��/Փ��1{npn�TYZ�d,1" ,��QL�����݈B�Ǭ+�º�1����:�hmo+E�����H��ծ+��!����-��+]D��|��������	ʖO�~���s��)��+�0n�ZQK����)B�	n�Y5�ۻO�C��
���a������N���=��wM|�G6I�9-���3��n�U>�9�d��0~�wS����u�H���=��tY/��@<M���]���|��F���#�䜷cn��'����q�����<�&w�g,W�;� �>=U�{F}�bj�0��3ą�r	��{X�ϋ�d!�. �n��i*�����y��d��,[�X����.��v�|
�����eU�������+P-�f�'_l'תVe�R�C�4��4 ���D��o=��]?���[�v�^�V�Y����=-e~�!A���3�����0�++�QT�뗰����׿V��x��mV��z[�7pY�g�hL� ����ʽ�7)�]$j�L
����x�E�H{�U�n�F �I���%��	�^L����٠D�:SG���X�qx.t�@�����65jj���+B�V:��Bm�EbF��2��踫�[��EI���u�!Oo�p�\최�f���>��vb�u�� e��g�t����N�_}�!73���³lE��<;�R�֚����F_�A+IV�\��o��(l�..���e?���J��}��D�{���C�~O�y�/�O�xf�b��>�[��#�:Y�MY�m��):�����ŭ�����/����'��@rj-����c_��>^�H�0�td���<�f�Ă�Ɠ(��F5�}�㑯��""��"�faq���r�ޢ�sA�X�}��Wt�)&�L�IL0˃1���Wa��-tZ|�x��gH��0�!b3��O���][n殰@�۞:�����n��T	������5��Q�_>��W���Cт�<9N`���.:�/c��걂��]�/=�f9��5�����������~�
��ߏ���N��3��"�'h�Β&Ah'�2C�
"�����([.������9@
�@%jk��lr}9޹�D�A�vl@Å��>��Ϛ7�LB*�����|��v0𾞝li,�q_-��������љ�y,|Ʉ�ޥt`M-�ȧ��E��X�������כ��e�K�)�(�:�6zG1+�J��f�oؐݢ�����x�� ���x_,��.܇�Qɢ2����_B��RխA�"*�]��+��KEG�V����V1�����|A��:I=�z��b���Xe&���v��\k]#��QѶQ�|k94��U�7	W/·�Mt����ʬ�?0yH{�r �h�U3\��c��30�Џ���L�;Ƌ�>�N5�E�q?��������A���$� �wЗ<m�c��CpaA��zqj��+���yFt���C�+ވ�k!<A��&�[JMj�.�SL��#��`���J^����bDA�>q������{�o�}�i��A���Qy��]� ��n�W�H^��]C�n.�M�f�=�W�F�ޚ]���&ytj~ ��R_j��#��o�>
Q����+j��.������ϵ�_����P�#΁���@���k��ȱF����D=��AZF\�~(p"~M�c�{��m�����ދdf���[�1�m����C9N��"Yn�.\���8���Ph���c�L%@:����2T�� �a �tq�ݎ�Fx��d�����pBjH�4Ն3B"�qt}TGj��"\������-a��r<�_��`�2+s&]��C�b�Y����.��~�����a3q�ߣD����E�$��Ρ<�?��j�T_H
LF#�۰�h�gf��mЈ"�l��C�E�0��%)�t����快�U̶��u�oW�:���zj&�ԾYtB��y���A:��2�-5q�3~�Pw`)z=_�hm<�����g�XՓȮA��|��ֲadw��vL�"�n��Gp�ʗ.�pM҈�\#d�]B��5��������(X91�#��ǲI���K���\ ?�h6�a��<><oNz�b\u�4��q6o�b� =�"U/���i6s`4e,�6��>�vv��0X/h</�b/sF.��ٌ�l�~xBlV��y����Y��13���pJ(�w�M�ep�):�!�z��	��ò�6�� g~8�UR��U5$z�3z�qf�J��<�~�t��ژ]�m��o</=1wbZe'Ϛ���a~c�\�3����mJ'c���S�o�N� ҎnPGG7�1��Pm�	��L�>Hm�.MQ���O]{�;D�v����F��?�e�#Q�pL�Yb��y{�ૅ�D䶖CUY�h�L�Q7RK��8�gJ�Y�tOj�%qOg�L�a���s9��^������i����8���u�%����H�7�ͺ�6?y��J�X�B.���3(!�Y	���Ga�d��!qw�ʌ��ǢLǇ+�N.�W 7H"�@�H��Trr+��Cf�B'-s��p����r�RB�����r����mr��s1��D�K磇9�h�Ht�( |���'����et�3^�J&m�V��;G6k8.��DYD��mC�wU�"��m�,���Ɉ�h����)��B�7��0�;��"����'�;�Bt'^��mĚ�r���(�/�X>�<RN���o�뉰H e�����a��t��� ��J��^%8ʫ��ɰ  �����9��Uf����m�y��U:�V�GtE�o;-����+��a^y�e�&�?x�c� 8�pq�����t��5:�%�Cj�3�[�3~y�Q4}:�TOv�uS��ꙒN�nu��9���'�ߔ�&/����=Ð��m�p&��K Q3<��{ۄ��	���Yo����:�jV_X���2��{`��H�����D}�1Y�a��q��Be4Ĥ�#x�.w�%�7���<�1~
&O��uWcw8LU�;��!ZK�P���)�����X�<=�:E�0�P��$�;��W��  �g;+�?�h_f����=y&���'rK�i����<��b4f�E`�Ի�n����T89&�'����t��-aG����X�"��ﮒ#@\�{��7H�"a�ğC�^�a%���3:�1>�[������t�z������g�k_t:@�2"gdof��8Z�~�p�.�W1�>�VY�q��x����H�W�a���0P%�d垱/w4���|���݉M��9�9�yT'd+h@�hU�x�F���5��j���^�NK����p)�/��\h�Iʒ��w{L.)��^2����Z'�W�8N%cK�3���sW7�{��9hqP/�o����Y5�"��6��=�OO��=�e���"S���h鰺��9WΝ�ĝhu@R����H`��)�_�G�#?�a�8����H�l�G�ز��3�P��z������q̠��pIuV�O��|BC�`�Ze�Q�z˷��B�H��FDp�d��O�7+y���؈|����R�9-����|&sc1;�5C�=l��D{{��ۦ�J2�-H���cj�-T��E���"��?���V	��7�H�
@�hc��d�B�n�kC�B~��,S��b%��Ψ��?N�Y�3E�)m�����gS#�\|t�������8�E�g�+@�K��kU�x�g��/��ڄ����2J#�I'��g
�Ga&� 7����;m
U&���G�@��!:S1S�2ɩ��� 3��S��u]��j׃��c+��4���q6[ڑ�{��_V9�!q�LbPr����i�m3�U���nȂ P���nB}�ziaeS<�|���4�A��y�L���)���:�;���d�)sb��H-�(L��ԇ���OƭgO�$S����Y}�V�"�
'c���kh������s@mC:2����_F�(9�K�>�[f��p��xݖ��5����9T%�����H=B¤+Ɯ��A.�޻��:h�y����.̢(3�N"(��b���3����3�v�rpl�����.#,�x��f���>M���IY,�*{���ķ�$����S��׶S�5d�#��r��̿�����B�D�@4�B�_�L+��m�Jݓ�
�����^�UJ�h	����F�rL����u�TszhEX����tC�z���Qf<�ط B�G�-��,c	̱�Kg�6��t0�T�6���z*�U J��� �F8��lmz�T�)���G�Jeȟ��*�M�q��N7-��Q8@��2�R�t��D'��v�|xl %�n���	~�d⋢�J�*.u�>@��J��X�YXVT3éx�.�����naI��͒�N�E],N��އ�ȥ�����O4ς�K�B��=��hhi�EGK���]*#�b�ϼ߯~�k�z���9B�:��h������9���=9�'[�e1$z؊��y'\�%��R:1�y48�Z��*p֗���^���8H����l��H���c��˙��ب�]���n�h�GO(����E�����O�c���ч|�q�^���&?��T2��Ҳ\�y(������R!2��&����a�4�	DA��iU�+=M�f]���&e�zᲊM�`��r�1$�"]@��,�WF�hd��Q�L�%ig��cf8>
�*�=��Gf��mA�R���DwX�JC���7n����}���������u��,��s?�����{D�j�^��WA��8��e�,�vQ�o��97^���J��	��eT�O%uOP�"N;9ĺ�
JGh?c�lBx�H����D�0��z�Zp��eJ��D�����+G3NE�-��1�/)�	��n�VxSa��L<f�;���$��,Ec~�����vq�^b�#��L�������_��RT�D�d6"�$�7q����"!������G	�B��ͽ�P�9< ���'@o�� e�(�_�U��˺�A����3\LB牒iF��C�_>���9�V�,��4`��O7��ߴ�j��^;Y�8�B3"ۥǊ���)}�$p<��*�6󥗂�wtP��ǧ�����)���{�"���S�2-�$�C����M�s�i�����i�Zo�C��7ƃ�����~��Ɩ�F����S�hF�k����OYu��DF���͉c;�7�T^��%��h���,��|cJXo�i�/�z��m��r�3��B6���"Q��eJ�Yn��8g���@�4�'���|�ڮ ���_��v�6�n���y�Ҧg/YM	`��S�c�-�|5g9LCc2O�`a�I�'5"�bto��N+����p�e@��zQgZ:�_Y�4���2�J�饓��&�ޢ�ԃ�1�@�t�'g�D�S�P[�5FoK��H�"*,�ݒB��i�o�ݟ���]֖$w'��.st�/G�m_�W�jȏE�����M�km���q���z�8�w6��[d�|j�&���+�x��6i ,�z�v��,�/{��tr�嵥�bO4��;R�d�tU~�=��:��b�`~��� �����L�
��RuQr�v}�i�7���f��+�S0'���N%���Dxp0���7����?��������v{�XU�oHb�:k�*|d���Xe��P,3 ��]\�q�����f���� 1�]G��

����Q�ʨt~jz��vmڒ�����q74�� ����y�k�����7��<�w+��]�$���g+����!ZD�I�'�l��oi٢�љ������ns<���=��9 W4ۮ���-���/���ﮄ���?շ��
%G��>�Q�ZK�y"ֳ�D�Qh�\�� �,~�}z�} ��v7����N�ܞ��^��-N�h��4���2D�,���i]���������iW�5N�X>L���<M�����L��!��&���o�K^MΩ���>�W![>��;	�O��`5����l��n�Q����'�L�As�T!�GY	Y)��l1�z?S���ɸ���U~�(�Y�X&��%֖��f7}͐�p[{��F����@N件���EL9{�X,�4X��M*��g\��.dl���"��6�s�`��>�#>�u�,&�t���J����XOy��hT�Ѯ�:Y�Z�ܺ��è������h�t�ɠ�w��{˵\�Lu6$>��^?���nu kR�~~���S�/�j��,��� �I`�����i�ڎY�[?6-w'��4��C�=���lJG�+���N��/G��7OW1`�����(MXE���1Z�BwC�y�� �ux�xl)2|b$\n�2J��f �L�@Ͳ�`vx���Z��T$%*��i��p�&�y�W�c��@~�Y�#�v�אꩿ�����]��K8Y��ǉ�;�b~�����.9� S0����C�sp��\��f�X���ݠ[�h�?9��4���d�>�j�����60A���h��aBS�3B��;C�@�#Ԧ�;��8�H��V�?��}�ך>eGXU _�g6v�F
}DO����4��J}�Mĺ2D��0�/���z3=L/`��Ӂ
������E�U0�ҭ?Qla�F�=}��;X���nD����4`{��:=�:t&0��4Q2���R֛g�Ң[�^z�`� ���9��Q5Xێ����U��1����+�����888�a���kZa&F��f���a�YAl<:^��A�S�h��FY��Gj��HE��X�R�@�]��T�E?�D��k��	G"�P�����8�'��D!�1�뿭M%��`��^���Vڈ�*esTUȹ7�e̲��w���Ў� �?��=V�d��!y���#���'!9��u�W����7}���"��;���b�zz��Uq��-��o9��"p�j�~^�f"�3�BIaz��"��.7���g�D�B����j6��}F>l���MZ�\����.e-�#��g��sH�|<��@�!:)��:���6��Ī>�!�1�u#��j0m�&-����g�����u�)(�g���c�?���L�hi���W���7nuWժl��3����*�`u�_	{k�"���|=K<�hO�ZȠ����36 �h7���T�"Pf�<��0�����w���(�ڼ#��z�v�h7�
gu�>�y�`���i<B&t��k���6WH��~�-��g�^>�fs넚n�Sސ�~��U���j ��䪦�|n|��JҧL%���V�����I��%��#�09Mҧx*⡿+�bphJ�7d���JkV]�wI��Y=��H炡Tqp2f��~�A4�?�q����s�1e"�Wn�C�٨?���T���?�!(��N��E�ޕ�){�-Z0�q�S�!�<T�����E�qȳS:-΋]�����̵6���(G�1��SHY���H�����3�~��a�w��s��Z[</������P��v���;ɻ�ҡ�ߺ�z��U�x�xa���mp�]�n��]�I�Oݛ�C�X�������Z_0� o�i`���]1?@�9Q�<;�;���:.�F��0h����F��D+� �z�~�~�鹤����Z�q���pTL�Q�yl��)���c8ꎻ�! �{#>q��{z�b�m��x+��2��Zt-ܖ0��H���"�MeTiS*�T����aۿ\��G=w&�/j�1@_��4���Mw�����]�~k%��C����!�OWe9-T=�(��q�,(�v.�K�p/T�Їa��<4>=�v$Z�t'������80��q���f�{���d��<��Р��PLm6����؆)���m�p�A��倪 	g_d8����;��,g~���N�S���bm��?��0gWH�p���<'��#��6Fz=��ygv��`8�hϯe�t?��6s��U��Z���pX*P8 ��7[|Ŋ��N� cזl"&��@��`[K�|�%��)}oG7V���T���ا�˭���3"��NW���C�c�B��������̙rK�6�l�� 0v��O���ek9�E-%��J{���Z�9� ��2=ʐ�W0Q�8
R�Ax�Y*���a1�ދM$�DN< *�]���ڒS��,��q����N<[���v]$�&r��LC0���kп;)�˝'�o%Q�8~�xb䝎 ?�u����6�I� �f��o4:��Y���l/1���v;Ƿ �}�"�u+�'�ҕ��nxN��N��IO���o So�1�l� p��7ɸ��J.m����#�ZZ��I#㮚�X��!I���'S�s�tƢL���[�e�=ع��LI
��|��ӑjE?τ��G��M.o���;�^�(C:鬶���V�࿃����?��^�*�H�T�Yo]�<���m|8@�9\�ڮs�
(��g���_5��ͳ-z�S�~�r�5���")��5���j����r?z���Ud1��d���u��7f�te.jB����{�,Z`�9�/J?�qN_=����n?��%�x�.�WDI�}��O�xw�/fhi[�:M�
%(�Q1��%�2���6�"�u{��J�O�O#Z�~^/�$_��N�G|��:K^�=;w̱�ƛ��gH
�0����vW`�t��u_'!��~a7�N���Kc[�L�8Y0�\R���#V^�� �5c+b���"q2��;�;�|��$�sQ*Kp�&�Wt���
�-�i֦���wY�W��1^�h�(IZt����:�������_r�nMُf�^QX�!V�]�V5yf�V�@�IxH����)�$5�or3�z�J��F��WV�X����ȗ2�Fu;�����U��p+�aO����nȪⓟ�b��v���?�������k��ԴO����|@�[����,��L��
#�Q�-�,5�7� 4|�#�=n�N�lʅǢ����Ɇ�=(魖A����Q���Dɶ"w�wS'��o{������~
�eF[�ʁ!�dٺ[�Bp(�}�_����}@�cN���q�y0�!��	I�t=J������0�k�����������q'u�t��7Q��iw�ۇ!�ȷp@@`w�>�Fds#f��d$�Hv_u���_$v#^X��W�W�?h���w\h[�C	������M�� �2�>��	�_}a�d�Yyڳ��r�pM��x�\�N&��9����@1�7k�'n^@�~�K���+uQkK���R����2[���y 9@W^�M/�Ty�I������f@�kOG��qG�<��'��l�Qa��S�v�E�����bjR>���Jpy$�8�W�BE������w�ܨƲ���UT:`������k���}!��4Y�%��l�YH
k�����U�`�ٕ�Wq�� ����ņ#}�J�4����e.(�ތ�]�*:�w*>��Uw‿'�%���1'�z#����M��&��V�}�j���'m;�
���׊ԶX�b��V�q�j�qB�[k��D�~���m�R�.�����ӈ` �R�Q~�bn~�'ө'!o�ؼkjo��Ƚ��L�yI&]�����5[#�ZTh"�M-��W��)JH�c���R����E`�/��^�<�ےxx�
=)4�fL:^�v���G�sQ .L��P�32�>�/��m�	��h}��]��f�eɉdz��Q��.�����tF�C��z�����4!F�̱1��v����3���`f$��R�a��IR��*�+��p����m��I�6��!eK�pW=�&/���.�y��HEN���nh8v�b	�qM�%�Az���X�����s`�'U�,���:4����3�gO*^�Ԅwʍ1,dP�j`="���\���Qx��b�I�	�Px 5�|��ڍϦ	����W��=�s#��&���	Uu{lu��~{�ũE,���q���ױ��S�47��)���{V7Mm���Z�`���;)�ȼ{|c��y"�im��T��٧2�ϓV"2v`�.��=";��p��:=�7�E-O,5o��3�!@c��ꄸ.�o����;����P�X)��?5��خa��T�9p�2T����88p��ǚ
��{dv�0�mɳ����uU��ڦ!�7��\�4�Jl���J�{��W9���>Ȑ��Vż�&!q���;���/It���"��Fx��@�u��'|8�%e���\R�>l��H�@~���j�i �+ �Ǯ��B��y�D�X5\�w%�q$,L�[z��v��s�ԕ�V���ʶ%�{~٬F���0T-�)w+C;:I�Q'�1�G�!o.-?�$>Iҕ��1�臈7�^���&�TM{��g�,_���_ Q�\1V揻R\���M#\�R�����*F��O_���7��!��\��S��f���(���[kڜҕ�����,�����u3P���7�O�W�C�h�͗��@�.?����T%�(=Z��d7S|z���Ԛ�Oex=��A*��ݨ��N�%ݐ���6���Ⱥ!�le�(��a��<�_��,�U2)zԺ�sjJ�oM���E�����ыC�s�)������v�ihM ��뽞�ݛ��0���;zZ�*�}������$@R�����3k�J�W����$S�`���^�hD�5Ub�$i�q�$�X��QS���Nw:F56ў��� �	8��N|��/�yu���|=%�`rn�89U��O:��L-���\5�*[T��� bF!�(�fc��lh��M#x�����k\����f|�sŒy��u��t�cv��6 �>�7V��e9;-d��(��0|A*ˎ\�מ}��O��j���L�iU���_v5>��?���H��/����A')�1����&�'r�t��`��t���Z�$�Y�I����t*�W_�� ռ%�4yGcY<��#��D=�Tc<e/L��'��?n�T��@���r�E��S^,�e��J�<D��-�.C �8��4�s5{g�G!O�y%��9�;��Si���|@"K���Ѐ���A#dE���6*n~$/���~x"��Υ6O|�`�C�E�@/Tq�ڥ�j�(�=�I�����w�������P��F�ޒ�Jj6N�����E�P�]f{Ę�Tޭ��cC|��������<�Q{(�S�9��UR���o�\L������*[��O]bDn]>���~�O_��%ٽc�C�`����N����eI8�ZqM�ٰ�&��|�ѻ���vt����J���˦R��޿~�0������ ��n��˧VTJ���:�5AxQ��%c���7'��8�!��VJp�>��4\���U��0h���d�%*���/���?֎���h������ە���<�ti+����R�Ґ][�$J?�x?bd��mU��!Jlr)&��B��/�nA�?�=���)-V���7���!Y2���o��!��Z�^ZH͵��-(-!Cq�RU�а��|d�K�@��[��Y�Ԙ^OѐII���f�⎯����ߐ@ʉ����ct�ĉzb�O�}@���G+�o��A��P�\�?�*�Xg�w��:_j� 8�:�������7x!��\�����u(�� ���FT�&߉����!�Q�<�_��:�cY,�~k�-�
�x�:�w@n �}cd����q��J���&ԓ�\��� �������خ5Q1  �HHo��^^��lԬ���8�]n��l�4~�����i����7���]�.;��`[�З�Q��F�M]�$�?�v���M_5�E����aV�R�F�}��)�v܍�Jr����g��x{���~����J������Y�e�h�PϰwsŞ�s�$����ؠ�=;Q���HӔǪ'l�Q"j�R9��ctQ�į׫ٶ��};�v��pS;�W�%8����:��H���+>+�����{U�w=,�c@�"U=�A�`�Q�E�P�����T��8�02��e�$�p�IԊل��B�㱩� \sM��=�K�-miKI��JD�[&�u�a�P,`�q�����	���*I���!�A%_�Q�;���Ē�ރ� ���u���=�,34�����藦C��;��j��)c�Ċ�X��w�L"L�A! �XBT0 m��?}Nɇ kuw�pE7�%�����٩�Tă�H�("_v�\�0�_=
�#J�z[�+�����n�߹�e�A���'��Kz���^П����8����)�s���w�mo�]�
<PsF�К�£ ��v����|��ё�m�3&e�0~�.������#nv���L{��+T{k|��S�Q�����$�'�&^x���n)�Xث�c���x���ưQs�i�(���fi ���%E��:�Y�{	=�"����Ⱦ�,CŞ( �o��b����z�R��;z���+E�n��o
Tf\ؗE;�h\�7,�R��.�G����d]*P%�I�8���+o&k[
�K�KY��\�ba���x}����k�D5&s*�p[tK_��o�ƑJ��?>�'X4R��I$�τ)��D�u-y�=~l�9�ۄd�no����X�IB�~24�4_���⾳�t�����w���m�RB\D�	
d"3���<��u�\�f1�j?��lh��X
���$wc���'�,
��RZ�:�6z#N����g����.[�;��`@GϴhX���E�BC���-�� ��Ó�ϩ1y'r��;Ie;{i1���Z@nu~�ߙЊ\����C0ig���T<P�?������$wV��a�N���/k��1�Ϥ;���{P�ͣ?Q��J����g9�9�kq�󯔡��U.�5�E��5�v��IT!1��h�w��x��U��ʄ�^s'�$DD�&��$��
��e�b���	FL/��s�r��!�1=�����3�������J�M�š�I���R[���͖��C�е�S��nG��L�����N�ŝ���R���u\0U�9��Kހp�G�{t�R�J��D��k>���[�8��g�r���6�u�1.v3�����%��G�`�N+d�+ �F8���>�(!/���&�4F=h�ffE�=�l	�iB}��a�G;X�2��<ji�*��W���y���M̀�>Uw��dd�ܥJ�s��i��_�2f,��>�`�usEauv�A�tڋ�UդĹ�i��ϟK+H��>%�*�u���U~6�6��"����+Î����q�1��Ჯ�m��[���n���� (E�H�߷�|z���U��0G-�W�q
���=�-�o�.B4,�Xk,:Q�Z,١��`���"@	��ec��aRd������fB!�( �T4}Ui���8���lW���yq�R�����8�^����У�1V���m�Z[����Uy�U������o���ץ�3)Ԍ��	`k�η=T1�_M����4�[��I@kl��Dc�-펷dW���^ss%����LG~����3C�i]����?MB��T��ѹ�7�-BP���O���e�F �|�f�6s����86��P���.?���:�[���xB �H,5jF1u���g2m⛑F74�ƒ6��� 	�tI:(i�����h���8�F�׳����D!��R��7��bK;�1��-�������������i�W�N�@n������0�S�~�s0RUޑR�k���` ��nO?�,{�:�Y �p��������A�L0����*^�&��f� �%�����h�5fR�|�)�ȟ=��k8�Xs�������172~��>�0ɳ�������+�x`� Ui ��Sf(q�}�4��j�ڇ�,#I�}ZT�`ڻ��7A��(�� ���o4,��#�O�_�l�J��sR�<���ܰE�#��-,A�Xh�\2��~��wA]i�=\
�~^[�醫$��Ը@;�T��*��:J=���nӄ��  <�D˴�ڋ�����T����p�}��ځk�
�8n�\�#���:EM��:Ո�����p ǹ$u@��Gm��Y$L���ܺ�M`�1�?6����n���������Q��4�LlV�m��p�Whb����h��q{u %,�q�����#
�|�l6+)� ��'�E&d��m.�<���m�A=�c��&���r��Ȉ��5[�'�ݮ�z.�'���YvءTs矔Z�����p���"Regq�pT�<󗖨��.�C�!=����7D,��RށA�*<����`�NV�ɜ/đ\v�,殾���uuh�[�����-t��q�h'��F�6��9r[���v�F"K:��tt �Br���j��X�,�o#H�<�
[ ���O���1�o�B��<��O�Ivw�U�G(�zT�?Q�N���<�Z��a˫s	 �f��I#&��ik��vf|I$i[Ѡ��\f*���4&L�Lۃ�w,($Ǫ�qTl�n�����;X�C*>�<���%zU)O{�J%5��3@��m8�KZZ���P4Ċ��{d^��*˕�w!�d5�R[���,�O�i�&4&���Z{r�-� :u'6���ț�D4���t�j�j���w�Ѩ�J/��W@<P��Mh����΅~��ڂd��,{�GO<Ε�pm��|#3rf�]{⪳}͑�����\�ƅ��b���wH.qwiK����ƺ��}z�:E�ֆ�k�q�7��*�#'L��3�����Q�F�_a��&ڝ�<�P�"���ꔝ�|*a�o�����4�k��G�LT�c^1~�h�A�pfBR�6�0p�Tѐ��^d�=*��5�j8�Rp`��*�K�1_w�)�nM�Eb��(�k]�RYMçԣ@\j2�X��2��*��ͷ0_ߤ�n}�'����R��Q���EZ�UQvY�[����
n�),�no�}zG5Añ^3Qp�!�wE�I5�u>Rv�����V\L��Xk�t�W.�����AԺ�����y@�k�k�oc󗼋��z������!�\W�����&����=ŝ�Q�-�c
t��_Ѷ`�I�Gv�'�� AYU�C���	1��#鈄h�O��猛)6??<�Tvm>w3��Nuƭx�b�yׅ��je��*��!�9���z�8w�HQ��}B�_��(���O��S�?v��D(�8w��x.L^<3�������yjXU�	>W�А]�Y u�g�~�Б�2�J~�|���՚w'@�\��v��1��.U��Os�5�j�Ԣ:gY���K��'��H�����=Ғ|�6{��=�'�+Oe�i�!aU�ʿ�E�R1�W4����2iz�]V�X[��NQM�^�RS㌘�a��@V����l�rW��a�x����g�c���v�+�mR�z�B�0"��`{,���Wm3+�}���ؕJ_t1�hZ;1������"
)���{P�눙`��G�5�ه�e�a�eF*[A��F!
v��c!�sY"�7'�H��F,�[@�*j2����o`�?S�4l�=*��-Կ������[W�^�a�B���kd�y���t8����� Ziq��tBxM��[�աϪ����3ɦs�#w�_��� 8;�~���7���?���A�����R���ƌ'~�>O������q������ג]���/�K5.��^A� ���������51� 69av%7�u�٠���W�Y�P����Ou^�������0f�I��Q�g�M Tz ;�-����1Z)�7c7`���)��~�� T h�&W�盬=QE�����7���F�a�QcW�G��?��F�΀�q�Y�F�涷I��.�� #�����U}7�OQ\���1	C��{�K6��#O���M�!�Tg>��ne�PU$�~xTr� ����e\��@{W�C�T��TkaJ�T[���A&ϻ���5X9=]n���<�zM��^6E��[�+�&�D��G/�9s��dew�"�6��8��W 'Ns֝YA�.?P-.q��|ɥ���9�v������}Ew|6��JجƦ�iHD��5�@���Nݝ�P���Yے��! ���sX��E\15:���m4�`���"��JtO���=A�sKeƚz�!�Ã�w�YYX}��
�L~��@a�s�Y�.2}S�=ʢh���n�GϠJS���b�-ɣ�f}��B4�*�y(���	�]<	Jg�+�l))�j�qJ8������G���|v���ʚ����q����,׉Cb����Chˊвj����x��E�=��G��δ�}T���㷭���,
5j���lx=
tY�W0E.]�Ǳ��e-T��c�9�؄���u�&n!�z�����h�c�;��h�r0��[ֱq�-��,Y^�lӞ�;A�4E�	B�����i�*Gi��Qk�g/�#�o�C��)�}�)ܡ��O ��o�E����S�n��Q-�����/�	��@7p��֠�(����+W��B�@�� 1��Exb�+�"ʞ�7Csշ m+�k�]�����ˤז��Z��$dʶh"lxxǕ\��&�wӰ�%�s/�w.j{�$��~�wD siq�m��t�dQ��h�) ȃ��楱���6����@�g��^���ӆF�C�^=��@ɇA<%��`�����G1�uT���S��A�a/��R�?SQ$������"rK$ZӃzg�G�HG�h���7����N47'��9��\֣��/p����f�o2>tRM�d��h> Nk��m�(�Z��AݫP�y�@���r]�>�/�]��{knN�1�*f�S]4������>0m�������A���1Y�d��ź�7��%������AS%��%��an�Jsˇ/+ɼ�����	�E���D���[�x�+�m�b2��*��:6�we��OL@�˜<��I�	�[	$� ���C3,����� e��t^rw`b
���H]�2cǦ�|�qS�9֯��"~&0�r�c�}w�"lDR�8c�En�t�x���sI��x���އ�8� ��<6I5kz<C���n
V��5�ek��J
��| fg�8?�r<�ǩCǲ>�TxZsx{а�j�"ha�C3fJ�U�Tb�V��X��n���Յ�/:F}�h�`>"�GgpPw�QM����.K�5���b��t�]�sM��μ���%{���eh&�ȼ_�X%v����`Z�7����*��E.��������E��вsQ����S���˲�����҆� ~���G?����2����$���B�����4���Gɖ4X��j�@:c��&��7�h�1t��Z��Ah���&.af�D�5z��b0�2O��
R�g��P��o�`�j��E�o<����s���/�H�_	��E:��l�HwL3��<&*�����-����a�"��SF���I�۞��LJ��S�I[������V����笹�֊C2&�C ����@�6�4��s`U��() ����v��_M��6��-#�t�M�<�@cG�%��7���f�v�9�#�ɥhBs�rmF2��y�%���CE������LF�TN���ȉ�
c)�ྯ�/��J5y�i���A/~���4o����������@�zF`e#z�1�t#�@���hG���V��Ա �+��GG�wӯX��H*O���H�3{A軡������hf�'���Cg�
g5�m+O�D9Zx�;eP�@����
^�(����n߯:fs�U:뻝����WG�;���!��ٌj���6ʾF�/Lb\��D��D"Ͱ�J.��`�#��o"��w�Uc"�]U$��ECZj:v��0Gm�B�\.%�N�Qlj˽��4���X�ۧ���yAt+OEs�ܡ1f�w�r��{I����@�4����*5� �[y�G���i��ֹ^��Xb@PWZ`�=&-}네�[� z�;�V�����jF�8�G�\���͡��lNc�Df������l^�H���,���m��,�P��f�,�Zt�d�a���L� ����Q;�UϞ�9�}�����8�� �[M%�������C�G^L���X���i/d���Ǔ
�ɻRp��¤���"��By�_��}��H0���%��]�O�CJ���@�P����¿��Àɿ��q�-�6`���F:v�x@C�b(A�f�zȓ5�b�!.�> ��>͇��Ѳ��
K�,���I���+2��t��I�]c��:�m�K�pXOC���nA�K,����q#F�P��"���@�s�2����yF�tb]	y8����lJY����m��"y�v!r�_�i�J;4�x@���`H�*���5G��&��3{k����qE�q�9���d�6�m��QG-1�?hc,����h�Jz��y�#���ˬ��zg�t��ZkWm��ᡀPC��T7	Z����\��A|���"Q�y��5���wÈD��`#����[�����=PCD:�J�f�D*�Z9
��p�/�1�4j���O������g�&H.\4]�L-R�V?S۸�`U�gk"�}��G9XS�B�����`��v��m�y��Z��w�$�@�M��+�j�_�����0�F� BKu�R�1J����r�	"�F�W�j�Q&z�D��?�rK�O��Ze��҂  u@*�������Z걇����<�Pbx+�Ѳ���\?18��=N �����������E�'�OE�bf��	i�C GeϚG�j��W���JfkL�0os�i�!�d�f�֫�����dq��L�����I�RN�0?@v��	T�p��`�����%�\'<��}+�}ݥ�� ]<C-� �d��ؔ/�
3T�!<2t!<4�����OTM���v�U�KMp��!�֑kf:�kb!IAEX�k�{�����A�j��� ����'=s��%-��>##���Z�P���n��7`PJ�"�����td�GRu�){@4Ī����!��mn�׮�R!���I�ߛ�v\mW��q�����Q9P��%����Q��a&ph�aO�;��G��� I�}9�r9S��Z6��}�[�t����斤;��P�!7r����L0�%p1��I���{�[FtH�(��I�_5\�p4�*��#PkF�֞c�!	�$�'M�o{p�b��.��� �e┞���&-"0��TP�ح~H{a����lL��|�V��9��5:����Lj��ߜf�D�����K��U
uG���p���I7���<������o;BI��
�Ij-u����o�!5��H)����NX:H3_O�!WR"�V���Kؽ���=�|*���k<����zN~&ڭ���3�&>�+5.�MZ8��	~ٻ2�����2b��J�Z(Q��]��':o:��� ߿�_C{?Tk���z>�����6�Q6h�&|<�����pq�Y�R��cz�vI͒������u�c^���F&�=�J�S�����g��h3��Cݮu��C���V������̘ά{f3���H�K7�p�Z���jt~����oM*T4�s=6'ޔ�L��M�R�'/��s��9.���ŤwVI"0La�O��I	����n�S�V�,�R2�}�0F�2蚔P\b�'��.��d��/�������f�}��A����;�$�����_���Yi�,T����ifK��2D�r1k��w1�4�b!,�C&�B�w����3)����=M"�{{��ce(����R�R��	?��r���e� ��?� d(n�i1$ޜ��.r�,�짙֯a�y$4��|������������b�9`8SԍN��V[�Z2x	�2T�b)���rc�$X�$z�g�e*QŢ��sQ��g�*Uo�p�,�e��]�p��A���hR���b
c�- �6�r8�� �B"En�g�V�{�����7����Y2�9[���m���:�w8�:���--��^�Ҏ�x�x���I�L�3	IV_A�!��]^�n�'y�o~/6<(��ň�i@���@Hɵu�;ߣ��u�[�$~���.�(CW}�i���܋4np/�Z8~�;j�2a�� ��7A��r��
,$�g|�l-!\'��'�m-�<�p����GEڢך�v�K/��M�~���D�e�b�g���}_���H��
x{�Q,�^q#����e�s���wN�E7�J��Hu�hJ��E[�z����V��|`��ұ$&����G�_�rB
���,�Y�Q+��&���#A���3�� E(Е��談IO�SӋ#\^�F�Y^���EF�g��=+��y�Hr�D�����g �'�Qap�L��o�ܛ�D���J?Yk���WN½�x4�;�+���ݢ#b���р&��5��E�@P��������IN:`ݨ��l�a�\nC�<{},^��6 C_��1�J��8�j������}F%hn{t�S����pRb�e-'yvۍ���[7y���"�	xdq���(Wi��`�N���Fpjϲ�G��(�<eȔ`�-1�1�h����#����ǳ����.���0����dU��#����ڲ-�ulR�xT:.@loAХ�33�F�߼�Xcx���������a�bQ��;�7g��+�7x�řd��b���4x�{��)�|��$��T��u�F���}�E �\�����۪-�o����sO]w[�Յ��XlUg� �}�>h�R��3���ڎ�Y@  ��<*�ZkM�T��U8�a��*Q�����;��|I�
х�S�<�6��9S��q�}wƼ����g��gi*7sG���d�n��wJ*ە��<���5$����J�������T�楻���1.��|�1�U�l=K���v4��]���b�o�Cگ�z�X'�U���Z��]3ݔ�o��}0.8w�TʛK���h�.�_�C����*�ޓjNǭ�uA�*�����S��p\
�z,�Ӣ���n���B��O��k�z-�h�
h�=q?�!���*($��r(GU1��)��Ǵ�J��*��&��Z�V�gX���d��]�N&�;e/	ǜh�ˣ&�!�1�1W3��f{}�җ��rGB�mU�v�(1~�>½t�fL������p�D䍷P_p�k�8q*��ߩ�X��ڹ��^�dҽ"��b��WÔ��uXQ�[������~>�P�[��3^����m����6N	V���<m��50O�?�z�D��n��u$�[���&��CE���;��S�0Ιd��SDJhsxT�p1]�$�l����t7��ΰ��X�-�#��� �>�)k �F���Z�0{��-Y����R����r}P4i� ?� ��=O����C���ŉ.�a�p���X��|�Ϲ̭�dY�S/�$������iW�mP"߬���&Ɍ��T��*��)I�2�6L80����
a���!��!)�iwA8�b���]����^�4j]�Q�����~���j�⮰&�#[��������GFaҶhK@a�U$f?dV�E2���.�S��(e� �
nñ߁�w}�r9�mE��Y��t�T]>����EgyH�<�ٹvȫ�;��	���g"�����I!0��}Ϝ:��︽��q���Ơ����=�&wP;:[nYul�X�m��S����6��^��KoĠI%���({.�?�L(X�Lq��E�Ξ��A�eؿ=��~���� {e"=*?�0D-{�Ҵ��t�(�������~��̨�ko���XV����7�#���<8bP2'�Hdֵ�q�bu�����F��;��* ��cټ �Q^	P<w�u@�9<�b���T�F�h?j	UV�p�M�Q1[pi�:�w����}G�&{,эO3��}���	c�Eg>�RА
��mH��N!�8�B���Ac���$�`��-K�eE��[jpn�0',�GŘ��tZ�2���@`Pk�WһK,OK [���[��:�Ƴ�|��� Z���W�I/#���u���d��Nz�TEe����!1���|�c�$���[�i�S�PpMg)�V�Fd�W��t��1J�w����ynvEJd)_���S=#�7��3��o+"���AXG4�!~pj³P�`;v뙐��^cｐ8|Uw�j�&���X?�� ΄	�-��G9�xz��M��[�ok�����<���DС *a�(�ʹl�����V��a�}�W��h�f�Ƌ��Nﰱ�0@��b�=��$���p>*K��Fm����K��A�6n#�҅ti�tIty�*�{,.N���R��Ln��z�Tl
{���6?ei���R-���xU�\�����`�����Xy�7<)1���3���i��P�30�ҧ	��-SxO*M����������Ih�л��e�`Q�iI���<N���S��q��Ҳ�h~`�y⛪2_sFyCL�^{��wt��%<�)w��w���>:��X���Y���R F[-f� �l�s�a���с��>�0�8��YJ����dӓǚ�0�2/]�D�������6��h�|l�.�m�Զ��Q7����)��Z��<%�h=}:|��������L \� m#/�ps�?��>�q�э��ځ�����Zf����	3{«��&�q�;g�7ԋ�I�8�b>�S��@�v�a.a&����`b��N�aWE+[���pXlI�Ja~&�JPv��D��s�� Vz�tK��^˔�w���3gz ���ͳJ?��M������?Sᥡ%fw��<�Vx���)m��I0�VPJÂ��G���u�;U�nJa>,ZN2�z�`a`�B�uOp��	=)eB;��*�"P&���=*x�2:<h����I�'�'� Pkͅ������]Ζ��'�ּ�l�Y8����y��E�Q��w�����m�" �#m ���Ƨ�V����DN5��T�;�r Ә|
Ё-��WT�_��
("H��m܀�S�Z���	4[�@�_v�#+�����t��H[���,a.�"!x��M��F<}d��%b˝��?�@�$^��;���Hkd�X�'XB��WU3!�b�%���j�O�K�� ��n�x����T�K��)[Z ��g�߹`��b1����+>U�˦�*� ������,���l��)�2K4RX1�H��a£�/
y�zi	���&���{/j!7w�j�tb ���ns3�������9l��ʋ��H8�c�lQ]ޔ���L�d!J�ʵ�l������|N�\C{��U`����q���~�V���/�Q�x�i���<���KZ"����|�]/=7.P��KS��j�JGZ�����m�H
.'��?P~�G#0���L�J���A�튐�OT�t��v�C;�.�dآ&�`�I�^?l��«���zl�Ð=|�8�K?򪬢�j�����H��^NO��D%7�g�E��@q�VB�)�]F�|m�������7��2�wp.C�>N}�/��8L����^����;Q��?������/�~N�ҹ�6!&;�Z�Y�!�ӥ�z�Ҋ=��6�G�b���Yup���#HZ���� ����B�E/πM�p�1��rr����]�}1	�8�r�A�e�w���_4eF���/��ү|A�e�,�����K2��e{��3��x��	�k�4�����b��1�0�r�{;����i��j�Ԙ�!G�֏kF�6R̲�t��؃��Os39�-+S��x, {��B �f+�XtWAϳu~�nB@�%Wf����@��*��;���^�I�'���(���s�CsB4k"�[�՞o��]�<��q����
J�Zָ܇C�:�Ⱕ檴�[������$�� T<��ٛޒ��S���s�i��!#�SԴ�!~��|�׳��Z��(�KC�7�?��`&�#␣�[g�$�o�R�� ��VJ���j�ã�LG��)��s|8�w�+�Eie02$��\��\i��:*��y�?��y������x+ϧp^��i���.�#�@�h�h�턅;���	wO�[����M�᥍���*��b�d
D��S.NF��^��۟-��13���_!���,'N�Zn����@V�!l�j#؟�3�1q��ݠ������KR�x�"X^hn�E��Κ�1�r~�*�М�;jZ���H�H`�ry����e�⊧�V�����a0̍�O����ɧu�U��yM�"�*�6b��7
Ƽ R� �H�#�7'�,?F�J�7G]x%�	���OUD�� ��f�/)�.9��h��/-N�a��6� uH7d�7�Ft"�&�ި��h����e��Z�ƀf�
_��xo ���,�ҽ���.`W?%eH#y������Z��		�E�||�F�Z�i�\�uC�[Y+4�y�����w<q�-�Z�F� �a��?��9j�6k��Iw�&�+cB�0vq��0�����S��/��_� Ԃ̎�o�jX�B��`W>\�|.�T���=f`\2R2�F;�o�ETFz�Ì�L
L^lu�Eךg�R|*0��֢I��q�t*��Q����*&�>�+\�=p�Mu˺�A��g?��=���-��Z6ù`��R��Y��(���y<�w���,����ט���,��*Jb�bN�|���P�^#vhb2����l#��WG��}�Cji��c�7'%��K<���[�[k�k=G��#�e'oJHs�@���ٜ�[��Y�߹�N��[q�\%g�IS�ϰ��	>�o��Y��-x��kF�A$��l_R8v��Ix6��в���k�]V$	�%����`K_��d<��!f�>�£�9ZTQX]����o��-�)�$�����5�)6�L�~��<�\&��l!5G����`��{Zgp�G��A�ťx��=���'#9c�kW���er�O���\�����O���g���u��7����&�ݨ�VveiT��7�Z�\�$��$"�oĹ��]�8*(I~���o?pl���)<�,mx�:C)������.�)7�5�mH˛�x�X���0��:��K2<q�"O�Æ���v��n�j<��g�J����1��g�}C�&$W�$�t�P)㞉�]��})�)��oƨR��.u�*9�^w�{[^��\vS���z���Q)�J�wC:�j@M4.���)3�G4=����>nkJ����)�ai[|]˄0���������v�P�� �	x�x�D8h��6q�O���@���'�qH�!�>n��8��4���<Ya�."�G�|�XZ����$�I�G~�w3neY�(��>���{��C�>ǡ�_;�`�;,�q���f�<��z�p#�N�~�q�Ƴ�u�eȧ��G�:�g�`u�)07���K�=���� >�}A��`r
#y�w�]�-'��G�@<������^�F�)����~����TSi[���W}�nŭӟO��`A�Y4�U�"��T�� 2��#����e=�l��J�i���>\'E ��M8�U�_�M��F�����k6I]�Q�vQ��r�[�@�k�s��$3F����x�U��ӳ=1����B�͕���.���DṜ�,���������hx���7RG\1y.�dcRB嵣8HOa $0Ӻ�4<�\[`:��h�K�7�ӎh�/*X��n��N�Y�Ϣ�4]u��Ӱ�a� *QR�G<�m�¦���X����=��y�"^?F5�j*��~䙔�oZ�7V��בX4g��Bˮ�r>�zkc���~�h�����$B2�L-f�ӌ���S{HI*(.z���=B� p�K���X��d\j�bţa�r<|'��/Ԕ2e�"�nq��1���Wp���
�������|#���V���EU��:�F>���(�A�*)��!���|�c���}�$�J�)#��0 ��z���'��*��T���U)��֝�����bv���ݻ �.�ݽ$̧��O`}:�3:R6j��뜻�΁V���T�p ��^�k�n���T2܁�N�*}�5������V�fԻ�Qz1��%2$�j}��^JA���tF=��H��]gE�~�ҝ
�M{k�!Mp=1��`0�_7���ɱ���u�-�Q}
LG�|�S�<�u���
&�;iy�љ����$��)�93�u�h����[1�BF�G���,4PL�F�"������<�2��J2Mk"�8}�yv}tG49�l
9v�=���A��sl��2ch,�8�l�����	p�x�xj�ܣ����&��SG��=�v���8 �Ը��fH���R��&�v����'R�P�$���f�fIFJ��9��^������M��K%.<�0��ݻ�������O
v�3�uK�yǽb}@HbH���v�L�����-D��n�a ����u�ꦜ�ߒ�F�����y����Juo��,s߸&o�J���ZM���.��E����O�J��i�/����J��
j=����-���G�5��œ�1/���p*".��_�qQA|��gܥb��Se�r��y3�	�6*�������!����L
�"�GjR3RV�9�����z�8�,;]g��L	~z(Y�Dy�)��{�Z$��T@B�\쟠1����>�^����G����ߔ;n���D�A��,|�%髤���ǧ7��;6����%JRp�ie��T�|&������W��t0[��
�W3k�ۧ�B����n��?쐕��M��ӫ��Y�WGZ����Zd�J��'Uo ��?�j�҄Q�R�9O}�h��g�f�o�&8�ĿpCEI0�����$��`v}]��z�A�{�㌞!wH)��1�,�]_SA�KS��?��ml�� <S;h��6���f�W� ���X�?�j5�3d��?�0	"7�ps�MC���:_-R_sl�gFUVn�&3���������B�vb�,��pC�������$�����̃��M<�y���L�����5Pr�`���z
�b��t�OP����Nf�����gf�'��@oP��Ab��kS��9Y����G�w��k[D^�S$8����n�`�&�KLA6�o�?j��'�]���V����2րDNE������w�a�XY4�a �dM�NA�K.RiIiLq�	ӌ�:�-$|�6���cV��W�7�f�#�UP���\R�-MA<�?��Q�U��7JS{�k`iv�H����5D���H̢*���N�N�Y$�D{p��=���l��~w�8�ͽ֕�_����d	�aS�Y�]#�6(��K��PѢ����'���y!J�+���o�����l2����J�`��4�����S\9e�4W�2���Ge�mx�+\U�[�u��r��l���y�0�\�H:9X�:u����ߢ׼��:gTsD�!Ĺ�&�KxPd�ğ�����C"x����,�Q#�����QD��<@�rI�e�ch%_��,�����Q}�p�5��k(��]�u��l��ĺ8�r���#��N��灥|m�k�>h�MR�$��w3��?T5���M�ծ�����IRF�7A<����-����~���mKr���Dt�c�F1vKyԧ�cq���q���To����D�uK'C_Y���&r�T�zI���юC"��Y�������nCDlf
9���G�Ґ%�� �<�B1TI�ԏ�L ���ڠ��fJ�(�	KNe�*Rh��b5V#ܫ62�h�����p�]1>�Qo�a����_�7�ݹٰN?����������l���A{��ծM����r��,��7�D��sg�M��XL�#��ด�C�� ,��K�R(��o*W����V��vz�� R�����ĸ�����6�R
��*D�:��&���#����{�O�;�|{��_t����)�ڡ��;Kpu��e�%ޣ�4aq��G��ґ��q��ޔd�0�C������e�~��By��5w�2�疻����oS��O�U�pT? ѕ8m>�TUb�^�e\b�/.dx�xW����3�%�� {G�_��G��d��>��z�Ő����N����O���;s��b�Ε9!ׄ��^ޏe"�st=\�:�����pb�"/���[#�h��F]/oo�>-� -uw|����aX^�9[mɭ��UWƷ���]�T�H��L����XF���%Jp>>�b��too��'T�]@T���6z�0�\Q�e�QsU˱�A#a�9� OY����q��r~��n�p�&8#!�7Ui��)X���ǐ�{��7�Y�w6"��3V�Op���=��}��	�1�X0�S��k�x0Ic��,�h�jI�O����N��p@'��¡,��<�/;©��L8h;�i�^V�Yү`<v�{|NP���r'w�ce�������g�"蠁����K72u��E(���2��k��A��\K"Օ!l*��o�G¿�W��*���d������X��,�ߧv+$�u�*,��Ǜ���U/,�L�~��Y.�lu��5�]�����(g��w}4�S'ҋD�]@!'J	f(�F^J����8�%��G`�2��Ԧ��2@򌦙�n��I�6�1��f�,��kG���
?����\��VTFN+$�Xy�A��4�L�O�Ѯ��� t*��P�����OJqـ�z=�z�z�^v����y�J�����(^�e~�!��#Hx����J��N^�����/�}" �s9�5�Cѻ���2y��o/h��QR�Q=�:��צ��X��n�Ѵ����[z�t�z��j3�U��Lc��x%���;�n=�5q\�`��:g�Q|QBvR��8�i�e(#�]�s,�[
;٥���\�Yu�L�{Ŵ�q5u�}Ճw:��v�˫�oKET��{�����h]�h����J1��� Q��������Fۂ�[O��MP�S�l۫,ª�L�@b ����cE+(*�Ƣ��G��((f�~<]�h��0'�O��M.��_9�{ZB@y�β�"���͜{3�]�l��K��҉�i��(T_Z&�"�.��vD2��
��b��N��H��f�m�==�}�������	��9p	�DE�-Mۄ�s�)8�)�Z28}�1�e�����<(�'uS��ѵ���yjRy�+ץY�+X��z������Jy��!�槔�nO�N���@��R��RZ���_����B�FI�b~�����,�����r����9�'�5��y�k+f�ǓȨ�����0�ߢ9��1���!����������J�T�����Y�w��a�_?m9�ȅQ�Z#!�&r� ��
�-��Һ��Z�p���d��(S��OajE�'BJ��i��T��M�X�y��"�ϔ�m�*\@&.�@���&J�yC ����a��9�q_W�o����n�8}'z��f/�]�3�'1_�A�s|�4Lu��&�go�J�刬�P�c���r�oN��]4c7���s��$�_�Jx���d�i���g	I�U�(�.�Է[(j��}{Vv�z��eR��sڄ�\����G�$�HN w��V\�k�Wh`�[����N3��6�l�;����������$��S*BB��be�K���3-�ȎJ��s�Eeu6K�?Ҥ;�3��_R�?�%͌��N�{��d��;�o:h���64�ѭ�/$���'�ȧPc<f�3l�ϣ�lP)��� 7�a�>�5��]J8�y0$P��/ּn����m$��#��=7pࣆzM�4Λ���C��+�4����0�ny�"�rQ��'/	�^��RxZ+�?a۶vo����D�����9�x�ֻۜp~��-�?-�� 5��;�տ؎�h��q*�|��N�2'��FL�F��2���E�ڻMHV��.����@��0"���<�Ԕή|F�gw\�x�#m4�5����C��Z^�d9�i�q��w����aL�³�V�û�rjTș�W7R����v�[��Oꟗ}�2�"�?�!r�Uv�5n|�I��\��Fi���pq��Fhe�l!�Q��s�AM��ѣdMy��K?��R4ȓ�V��o(9��S&R�#{qw�ׇP�y�Ș���
w��ۍ ���d��CM�m���'!�,gBb��+�/uK;�>�'0��v�q�͇a.�bx�w�a��~$���0y�Ub��jY�˥�,]����)�]Sd���I�]����8
v-��%�7��jߊ���J����a;����(*����q�pV�	��V��E���Xh�#Z�5*z^�#��j(j��?w�-��}t�~�O'� �:p��m�H�B�A�����O�_]���[������$�b��C�s�;c�a�Ղ�Dΐh�]h/�a`ў�˻�_ҔQO��M/Dh�P���1�8�KAL��X]���<01�|.����xjlQFD����B�DYC��ت?���4^Zj���oF��������]��7�q�O���Sў͈Ro,�d�h�<�Sť����n�Zk����n���l�(l�����5�\�"�Z��\8�aC����qs��YF 1�[��C�f)�X<DڍE_�j4|����#�?y�[p����b�b��3{��c�����I�U6�.��r�@��f��Gc��J�n���}�@����/>���O�������x��<��h��2ƓK��}xac����?h}�F;1z�L�a���;z��65���/�_�p�N���/|�Z3�$��gNdO;�
.��6"�5���#x/����|�k�,��r����4�B�ԍj�v�
I��
x�8=�˱�ǁTDMQ��'x �z���G]�z����~������cA��QNB��U�+�wh����!���抓�i��m�܊V����U�侤��M6��.,�4|f7�>��c!��q" ZÉ�0� L�g(ݧ3�l�P�c�AX��&���:I'S�(}U!�Q�����(�e�s<�l���%(|�@��ny-vէh����f�$�y���Y���'�_Pc
�4!x�!ZvG�S��oV3�n}X�,g��A��@k�s�`Z����p�k��Ӛ��b8-���Ǳ	�t�����b?@�#�e�eiR�h��o�H��=�=O/~�J6��*g�?u�f2�k�4̴�mڄ�*R1�=�`A��۽�b;P�d�G�R\�t؜����S=����u���t[���/���m�e�)�����Z�MʍZ�b�3 ��v�ME�x4�0G�X��^1����#
]3ߴ�(� ���G��{~���A��E}���+���E����:��-�jq[��)㏗㗰.Y�����=qE��:&ρ2����P�p�5�̶���;Gd���F�CU�����V& �`�	��$����G�+���{�c/ל|���,)�ޖ���#�ʭ���� &Tz���(V��)M��xt`��=,,�����C�ͬ���K�m��%,E�$|SA��CO�U�]����4��sI���
� �Dx㦌�j6��Ӗ�\_��A+�����qK�~�Í��x𕚮�H��YᏳ�<��Q���F0�=�&d�AۜƠ8����;���:��P�Xm��030�&�#�T�8��Q��ڟ?x�	�e�=vT90Yе�~r�S����PDR����9D@ R �yew �y�\�#Y�^?��WJ���I����r*ӣz�Ht��ȭ�Y[ݰ�f+�*yPt��I����f����"��QhR���ʦQYB�i���$=�1za{�B����TL{e��� k�����Q�%ݒT���M8�!tw�Q���ZWE#{�>׳N�ߓb��R���X�$��)���:@us��O�����Ѻ{Ah�i��������<�B'3A�*�:�����V?"uE`qm̿�Ԓ{�h���}YW;K��륗}�`�����ɩ��w��*��w�E�s�̠��`63V� ����dd�Yj�md,��u����
��6��sqʛ�6�c��p�l���/���P �7.2=#5����<��S�=(��O?�<���`��#g��t���Nt�Ι�Ӷ)E�K�:�^V�)OXPS��ե=��r��#�<��Vh[8�=sk��ߗ�ŏ�;�6���1�5�oX<�l�򞦻ISo��%�=�+7C�[�L��m�U�����>$��
HOԏ��`wpӴ6���E��F��l��i�eL��W�����;3����5O2�X���lw��Ч�1i����B�woT5�;N���Q�<{��F����D礞}���G`L,kC�1wǽ�<=�:�:�d���R�l�7 ��Sx�|E���T�4�������:�H��k�B�|���Լ(.fCt��5
��������u�Ȑ��Ԩ�L*��r��X�U�>�uF!T�ɲ�Pt��.�O�S�7F�Z(B�*'�EZij��?8C�"@=>@L&� �QE�q�`})��d�R?�푑��o�d;s�r�h9m�f�h���r�'W�
K����N�]�E��PUJl=?�`^�x�+</��S�����������h9��m0ͻ�/x��KRP��	�wg=�L�j��YQ!���X�{�Nf�a� <`Q�8��
��A��V!^�����T���uw\�c��m`lUU;|��K8 ��g{���g&I�;��;�)���[�3�<B��SI��
�/�Ꞡ�$�cx֔�g�b�z����U���9RY=N�F٫dvGZȡKT?�b�Yje+���y��]	�_�=�:K�c�}���խ�_�_�g��Hg�D��`�t24Z��&�( 8�A�鋫(�sKבD��R�+;���P��9E�K������Lv'ZM'�u����&j-ᦚ���o4��s�t�2���&ώ[j�-�G��j�㇑[u!L3���y�Y7�b�7����y����CNߵ�}/X#�{X[ω�T��we������㍐��Dңe�8�����v�?���[:�8Ӗ�;u9���i�B�b҇�x��TH�tJq���} $U�+��`/3���`�����-
Y)	F�&�aX��4EWϊPy��N�Bx����ʚ����Vx��B^o�ք�u`a��v��:�Æ�x��u$lG.�]�V26�����
�� *���hD��Q�g+qXKIk�\�5�a���s�)�K���0a�b�q.9Ewq��=3����4�1�����C֣�*�;��П��2w�x�BG�:Z︒�H���	af�r2`��G�m�nDsJ�t��.n��rf~�<��"�/��pz��`
�T��q~m��쾁Mެa�b�eN4M�s�s�I��w�g=p��'��T3�A�hY�%�	�8�B�Hp��$�JT�:ͪn�M ��}�T���b"�5Y����UNcE�J2�
 �E'�O-ɁxR��!��b��n�R#���T@��ܚO��k�V�����j�.5�ϖ	��Z�E�E�k���m_�̎�i���L���(�6ךڣ�@μz�԰��b�Z�q%;Ԁ@�N
c��Q�C����F�XAz���w)��(�NW�d�lY�#o=b�9NE��SŻc[��n�vீhj}��o<�W��K����G�������*�lO�0=a��>XX���gQ_�J䱫���GM2�s.�)�n�E��`'o�ӧ���#��Ĭ�H�ߝB�M���_~E��+T_n
����l�4>��U.a��^��^2�顮���c�sͶ�����P��`X�:�2@~�,���Q1zU)���-��J���VZ�zP�7��9�`�3r�����dI�s�s��w\X` X�>ڇ%T��.���PL�J�p�9�e3&!'�:V��4v}���?�� %,A��.�	t6�7�N_?w߿A��-�\y�w,��9��Iq������u�q�jp�۬k��'��c�-�-wz�j�8�GƖ/q�����̷�H�*�kq����6��sz�c.���E���Xl��󝏒�8Fw�my�O��(���žM +��n�C�K�E{9I�(p�����^�uڙ��4��ԍ��B��+ �_�M���sJ�?�]�/���jӜd ��yV�j�z�v^�*��c�+��n 9��&69���ݿ3y:��ŹZ���_zҀM9O%)K�xǊ'S�0�l���;���ѵ@�g>4�:`*w �+��'q	t�����3
�W����HV/f���(�z"!�~m.�j� �(��o��^�w}�KaL�U�D��M��X|���������5��B������T��|�L���S,Y�@\��Ş��7@�m^5=]C��Ě���D~+[fD�=e�v�gD����'��T ?�|�����a�u�NW�����҄I;ڦW	)��|"� �g�Y@�B(�WRK�۪Ye�������$�;�����!7Sm�	��93�I�+*|˽�}\�ǎN�r�t7E.V�j"�>�\� *����
O��t_��w!������^��D�����\K*H>2I��j�<z)��M�8������$"���1<�N�/ÈjG�t�;-^����qF&hl6���Vc(��Rr�a��3E%&cC$tP���D&cײ����80�42|1���� R�uZ��O$uz���*����!��/˚�bQ\8����gqҌ�ieD��({f� ������l��y�R����@��$s侄��)�5�P�aA�ʻ�8O���g��<Y��=S����g��/��4�ms�|)�Q�L�$�b�Yd���"��a�	xՂ�՜��͝�J��l}Qc"%H�܉�ג�K_�z��;�nH�������$�}pa8�����φe���ƟdD�L�6[��w7��Hԕm�h2���/�<�:���M�,x����Y�i�Ҭ*����f��F�EjJ���싵���!6���E
������n���陏:�� l,G��<R #|7�ًz7�4e����L؅�@bhY���<��}��oΠ7�W!�}���-�@�s�g����_ap���Y����02��b=X����hԍr�dM]���	��_�����aT1 ���v�ڢ�2Rs �mcLB����c�����utg~$5�����[����
�a���A'���,r����h����������SfZF�D:�t`V�H��#[��$���= 6����]ChW:�ĽFt�>�ăMT�:�zrB^��H�l��,��7bZ�����G�$4)1��(Y��?�AZo��zШJ˪�LA��Y�����J.t�$4���y �poJ���*�ˠ��DӋ��_�(�]�j���]�1��~1�#�)脛L�����ʌ8j�mT�(Qn��Գ=b��$՞k-��~a�0g\Z-kU����,U�������څc��?�1]M��YM�@~9F��T��p��TfP��[��$�F32r;Ծ�ϛ*���x���+��݌.�s�1�׉8+^�s?���s�YX�Ǥ�eo�b�� ����ϤF`�P5PZKuNjf[� u���_�O��É�_n�7�ۚ���o��p��(�βF�!{J�Flw����T��/෪��#��F��Y�L�cH��v`�]�HQh��pA���ܝ��7�;q~�ZRb:8d�ҁ��'�L���M qq��ք�{��B��Їq,�BU�P�L����Ij�עV�:v^trO�/c��Ti�睉�_�r:1]�3�J)��nr�\�j綰��8&�F�gY[z� � ?ۃ�$���_6;s��ҕ� �,��5�硵�'�=���,,����j��ŉ���d̼�������d��t��e�3��3�b*H;o�@���)߁���ll� 6��R���(�t���f ^�	�FU\��o+, �0l�60@�L%kNY����e6BU�s8���J�*�/ψ@1|FZ;�bF�����?�2D����hFĬ"p��ܛ�7s��@�����I�`��0@A����Z�0�$�Ȫ&=��v�+�k�틜���g[mdl�%	S����
q3Iox�9�p�����l�8C����r�%ޜ�M��~9�`��MB5l�n%~�(?���ť[�ғ-a9��E�8���V����o�����}~̉Hdm`��Q�|����(	mZ(w\UE
��Xdw��M�7/��R-����� �q���L�*��v& -���R�^h�{� ���B���k�D��aG�]��#�u���L��|	6�;ױ�vu��5'���ظ=��J�ES��|4��ã8��-������Z��8�ӱv��q��Fa�<���s�E��ZI�=�w؇Z��1ڄͤSZiL >���ԡ@�"��X�����7#�'g��Ϥ��� ��t�ѐ�=�k\��5]G����Y���:�MW�փ�>%�8�y�B��/[-B�{짋����mE1���l�8g?���sr���t�2f0�8���
�&��������  m�-�A)H3�w7���p�_���}��R�����3N���92���t][3L�G!�Z{l�<��-z�4����Ī��j�ދ �߷�2j&���,�o.�̆)Hp�u���P���6���Q�;i���}��y�2jk�Aό�b�~j�K�m�<�yy��H)�qNt$�!/������(�!������L�����_g�#�Υ(x-=dX��D��|�9a��q��0޿qǃX�p�a��C�/c���JR�P���F�/�V)�ZNM6=�����(���I�_5�k�RrZ	�9�D2K{%r�IQ�Wnt�8f��W;6�ny�mM@�K�&��F⟆�E��r��~���sN���RG��r`�"�mg;��$�]��a�t6�+�kbZ<��C]�߫q�zڬ1tV�/󗬸��G�8}{7�,:�"�;h%4��:�5��,�2[�0fM?m��9��P܁����.aVG�8����Η� }�}-��^��0u4����;���ί���?�PK���_dpV=�x���"�M�+NH�[P	|"��� ����a}tޤ!r��B�+�IT�Z���2j���%�CQ�X�Hm׌�o�ci��}<��j�F@\��d����\�9�=(���С5�O%*(�43�I�#���.{�]C��qF-�#�e���)�"�z�Lz�p�.�63��G�t	*$)��[ߗA4��Z0_us+�kX%��ڤ�U{���.nf�s�������h!qBt
�b֎�A��G%�Z!��o"Q��s�{'U_�������N�wҞ�rn�>�V��S�e�� qGL� � 2�����q���!��
�2'����8��2͉���	f\%8�P)���T��̩��[�^0�?|BV��zöL0����T�_�D";�*x,���G�W+T����R;J`�k���-��2� ��O$�C�e2��U�'t�/��'�O}��AI8d���'�ɟp�~�$X3�#��ú/7a���B>R�aN�K�|��n��V�qg�g*�a�eƶ��|�����NL���@ �R�e�JU�Ͽ*q*���=�K�z&&Ӽ7�	Q����}m��TO%;�L[��!���W:3/[�.zϠL�����K��ߴ�IX�Qcn/?v���R����ۀ�@A�W^t����=V,�؈=��$i�ö~�ݥB��ҋy�q�h;u1'� 9�+\=q�N��Wd�1�7�K�ƄSuj���S�I����pت�����	�����9�biGI��$�����<���������ч�Y�"���'F�H2���W/]�Z�(SiՉI��H��mY�fe�A1I���%bl.6��۽r"��t4i(K����:>pq�_�j<�4�����l�R��z�)���Sy:�[�D��4A�}����9¬!Kׇ���T�oA���iY�#�4h���ק�L��W�G�/��0��u������N�2 Gm��Q��JL�6~��*N�Q�Y��&t�;�K�#9\vv�y����X�xB��a	L̞oZ�Zo�|�ɥt����
�ެ��M�q[��Cw�Cў�Z��**�?�����AsG���7�6�2�ߙ3�W���5.Gh���jT�,_x3$�����,��e��i�m�?�w�P�֌�]}�8�7�9ϕbLJ�Hlmh ���<+����/7�#�ó�ys�GEм ��̧����NB͋��Ua$c�ִ� )�N�)���y�w$��Y��v��H��P�Q�HR�F��V��?d�h��g�b�Bb�����@�`�J�AE��P�֒���*+s<���]��|��<�Q|v2 �!{:p�}�Uh�@���q������a0�K)[W�Q1\���nJ 	w�N\)�M����UB6��������x�Nc��m�6�=̕�w/HƦ�)��NG: bB�~�u|�d��O`��";i9i$��]��m{���`c�3�i�FTS~˥N$G���;!F�*8���ꅏ�x���.9�G �g��@�X����41ϯ<�V��4�j�n��w�ۉ���~���\(�Bl�u
������)��Y0:UimfԌxW:R���}���p�F�&���<xj>�|Ҹ̗�K[��]lv�4$�Y�i��ݔy-�s_�[D�L	�'��o{M:9��g}�O�8P�C�Ҵ8<mΆaI.K߅[�F�Yt,U��M��c�I����2 �$���ErdA�$o�8U���#w��>�s�GyET���pF���(��RШ\�{�lC���anRc��/�9n8t�G��BT���I�S��x�w�w�@�
B�S!� ����5H���o�ǡ��Q��_'�gHĆ��揦��K�D�]�������O)Afl��� �
���;b�ot��cx�Y����F���=��7�I�!hay�I�o��������t���J���o�o�����0�9�s��u�C%6^s(���\r�SMqnZ�1��w�^P�s�E��o��Ù�3��E�Z(�U��|�=�#�]f-��I��P���ͼ<��Rcц� ��B�t�ӓfY�9�~1)_���
��
�
��EY�$=���&��z�����F9��uy����rH�\��<�ME��~��;�>3����*O�Md���$�����d��%H�{�� �J�5��	�lw�� �/e�9�4�)��YeGiÑ��^jbs8��
����C�2�K�7��'�r��g�/��°��0�0�eR;%�r3LE�#����^{<w2d8(D:=Dv�}���K�p�8����H�s�N�=M+�. ��vD�`��!��5Ӝ@B���z��7���7��d=W�[7�w��@c�(���o]��=Щ�:�ْ7�3�փ�<�:��F�{��H�C^6��;e{�A�j��y\kM�`#�}��j$ ��P�}���g����k �ב�|I���(�ޛ���M���qE��c��7l�H�N�A����C(�|@`�v��"�B4��H�ۦ�˴6��/�t���$;��6-ۍ{r9ڤc�Nqa��5mU��p9������7����H;����?�g�a��	W@&s�������b��M�*�V�"�S`}����Ю�n "��;	4�f
�-�����u�u+���:��~��~�&�d#1⓽��$aA�-H��)�7m���#���r$�GLT^�jv���Mi���SYU����Y�)��1v-�
����$�0v;rsX=p-Y2Ā �n�W$�㘳�Vi�&�n=��D���n� �uk�ĈY� 9(�Y� "?t����d%<cS�b���!OiZ����(�P�a�%8I���A����J�E�M�g�� ���>!JƝ�f�u�ٱ4�@��G��:`Q߶ 7��e�p� �Ǎ[S�ª	�]~S�f�	�|l\�� �]u��=���6������Y�_�TF���"#�G���,mհǀ�l*1��P�L."QF~wR�vk$F��a��.�[m,R��M�	�ERN�H!�w��/Ɗ=׽ޱ��u��ށ�F��DӖ�[)��j��Pk�
�j���=�Ѣ��i/z���� �����kv��i�k�U�fIE����x����my�w2�z?�hZ3lR�p<��U�7��QKv.\���b���'a�\��������畷=�H]Gut���7�f�we������ �9�Ml�M50�j�B>BBy�H�aS�[�5��_��`��/0˵���>���mt=���'oP���W��n�O�n�!�����ڴ���5��rBk��L�!��v�;H숝��\�wS2�9N)p��%��D�p��߸���V�@2C��j��,:�B�R{x(�-l1��n̓[J���e�����A�u[Z�Bbm�^��՘��\S�B�q:���B$l�,��e��GW�*M�,z٩7��<;�㚊1�9u��\����J`'1�7['4qS�$�b�QFe��ߝ;����1L%8H����wP�=TI��!b���`��w�H�"����z������O�D"Ĵ��_�� ��n"�0�b�aE�/u|3FO�Mh���"��Jv��=�1�$�L�L�����U�<�7Q��U(k��T���Qؗt6��R)#���OQ9��I�����ZQ{�en�C��5���K��$�[ſ�C��XY�'�7AɌ���:O�PK��'|ș�<]���$)��=~Z�5�_
;�*���Ʃ�J�!�?�_�Rۜb��O*�5�Ȟ��_p>N��?��Vi+ ���z�Id���9Ayʩq�*h)Csė�\!�~�G}����M��1�n|�^�8�\�+�h̢q70���Fr0��J�������sF���(�ZG!t-�)�8��	r�dO���n�9	H�v�'Emh��rX�O�	��;勲X��o�2]�s�����0���4�ډM�M	����8�<#���u]<�<�U�/��dm���Gp.H�qˡs��ݢğ�����e�����h&8��Ӯ�r��
c��uc���d��в�j�wsr�'p~�g�����(wM���'�Il��t̝���3F�Aۤ!��2��yfT�i#���,��=�8D�ܴ���Ȃ�*� I�ؖ����`)��Bӡggq�t֨Y��AW���d�M� :��h��K�VsaZ�̴�/���ˉ�yR�F��<<2�Qen�^|ȋFZ�����޲03�c&�2A�B�NA�O�U�(Qњ��Ӧ�y�Ʊ<gi3<�ev�DBRr���� �h�((O��I�>$8NX�˜QPc�|%ǀ�H%�?$;٬u��)+r��M�.����)YE�2�^T(����z�QŜ~R{d>DP;�A�.�!��������P�n�������ҿr�0�(�_�e�9~�=���(�zÂ-b>��|j=���,���X�L-�BXr�n�쓓K�N�VWQP��AMҲ.��-�g�ZmTo>^�h;�i{��4R�H���fa���O{^���|�1~�7�<�x������!�٩!Z�`���.b�!���֬�c�0�H���%�^��`"��P��%Û�rh(!�kDv�F��j��&��Lw���.���'&���螼�A3g�OS�n���������_���5�:2����-?�q8_��ȯ�A��D$�5}TR~��Rq����B�Щ���d`V�Px�J�$}S�(��10#���zb�s%���E�U�]@f��c��M�W�AB[4V$>!)��\��/��$������% g�)<ʭd;9��~n3�@��"�uG�7�f�}�:X5��0�^Ivb,j\!���K������S��̮��{DW��n�96��k^��ĝq[�V��]��s���-9W�$?LXh.Ú�2�r;o�Л�>�y_�k3"�Z=��M�2�]�N��"���|������}��L0V�^�ʉ_~�K�u����=uk�LS� ���\b7U&u��銹p���D����菤�����f��o V��F��I�8޾])�2o��i-r_9��p���$	n� ?$;&��q$���	3	+G�O��S���kׁ��+HjU�b��_��x���c�6f!B�I�dM?�ߪH:��y0���÷�X$���vb����P^q�j�@O/�b�9[���~�~yΎ&�yFf�{��G�B.k���vC�� �_��]Fʋ�V���[��\rM��h�
,@��j6�^�%����)h��<e�W��[��` �b9���Ү���9�'�d��:IHv��c�?C�n��&�|�q�p��u38KRj��@e,�s�e;Ű�{�z�b���ȗ����O���I5[�p`�s@oܜ�7�5^����eo7���f�����.����É�������>R;q���R�~=�9�o��`֠;�A�
��$V(7 \sz�]��ÒZ�vԊ���_X���S>�'Ǵ`$,
fؐ�/���ݸ�A�`~R$�����h���p���<����O������N����e���1b$�ű�t��9!h��"S�k����w��<k����
����}}6�{�#-z{l蜠�� �S\&��t���?���[^�9�Ie��!{P&�R���S^��e����m�6���V	��6��0	uℑ5���|t/�Lk��`���&e��ֈ��(QuQݤ�#�����ub���|=Hf2�Q�jjkxx��&\�`s��tk�&��}���~��8`׫��5	� +��-����j��᳖>����&����������'��s��J����݇��Z芾�{�Ǚ�n�8���
�9�ih�d���*�[	�p�W���	�JQڏ�<P���F�����[�,������Y�����95`�2M&5��Ǩ'[�3���F:zż��\�.D��������tڵF��o$8��O�b0]���SE��K9%0S������S�Ax�u
\�׆/��Y�����,2��$�A����xs[zz�l5��0x��!��ȯ���6]���d�s-�_L�U��A6��ee�C$��� ���S�z\��x}�TB���d�s�-�4 D�D��&ޟ�+MoG	�OY�e����pECE5�B���ӣ-.�ذ9��$n�F��6���4F+K��y��:�������8f!@lt��ݵ�E��e;�W��H3Xw��~n�Q�+V�	d%��ü����	�ȡLyt�)`Y��}�\�;m	gv��P�z��PVÓrL:��F;J����2VG9� 0Tj�|p~�V�xxA�dd���E-��	����]�`�I���](���_I0�$jn�PLo$GW��:�V��,���g��?��H�k�"LɴA#ӄ�k��(ш�C�=3���c�]�1���<^��;u�q�Pp�ڸ]�4$�i	Z4�l2�$󚮨>6��={0,�VǍB�3QF_���: �0k�`�ޡJ�j���$���(K`��Rmt@�=�:] �qb�͊��Px�HyϹ6���^8�3�'��{.s	N��ݍ��޹�/�����2�����G�x�v/$���Hj����e��r?�T9t�à%�K���mg�C��w�Iq&�hm/�����Z�E?s.&��<X��_�03k�8_���]���	�o�b|6�n \P9��pi�gY�ۂA6�=ŀ�..��ƉAX� �XI�ydg,�n�Q�GiF���(��j�x�%�1o1������F3w;�V�]�@_˗��ǐ��ک>�Vp����q���(}�%�@F�a���'<Ϥ���s0�X[�C��n�����7���H��-�t��/�g	�Kk�mԛ.�:�m�aR&����D��2�����7�{H�����t��$��PNI-�o&�u�<.�]І¡���C_������5�+�O���IZ��ވ�Hg�%��t��~Hb�=�QXZ���[.?q(�OA�}J:
�{��rOc������=8� |�*�z4�\"�Q �������8Ic���r���9^�ڶ�� 6z��U�ғb3�~��=`�bjS��9}�ϧ�S�V�N>i��T[���x\������������O�B׏�:�^N�Kgm����b���nꍉpB���S�(u)_T�v�y_��?�|0F�y	~���sP*��'�-Ay�(ENǹBcm˽i���1q�P��ϕ�R`<�`�����Q��oƀ�rM���R�-��T�*2�������孎�|qM<O�1a%&Į�.n^�E}�iȟYR&EB~+���΍c���z?�o��pU�#"\�SPn�{��2g��f�,"�JNf�|���J/����J�J&,̢e��R�6�O> 1��X��<�R�%�E�RV�C��+5P��k�^�N��n��L�_H� U(2f$5�R{��5i @Ѧ�>���E�[���".������0D��u�^t�D��3Zc��X�k`:�2��/�;����Ay�2���mA*@�4n]�p�Ȓ��_7��1&�>����wޟ��s�~��6@e4*�YJ� >5��w��cb����c��`��^4A{�n�.��&f*��i�y���_��T����lT�x�/m�+Ax�
�U#�~����D�w� �#�`=�
3 *B0͠7W@����u�p���(F�V��L�uג���(���2� ɪ�o
���p��{���`7��h�>7�D��+W���.?r�K�����u����w�$���?e�[����o�C\u��Hckj�U�=��V ZI���	"��>�V�vi���6x!�.6cQ��[U\*��B�I����~2%#��Fw�;�gs펢�Gi=���Q6�+h'����$rA�￑Y���Q�u@f5��W?K�r���޺>Nܔ�\_�}�G݇�G;�ǆ��V�A�_]QNŏՐ��)����Ȣ!]	^�_��U��Œ����6�ߤf�P{Y�)Eo�{���*W���2r��?�"L����j4f��R���h?�ɴ��a��E2B�y�c��' �L���:1�=b��W�E37��+��S����;N��0� �9�2�Z��w!�ṹ.tս��0�֎�6�z�_p+q���F�����=��%�Gs-,�uS������=��jeڊ���m#�R�ŒNɒ��ᒗ(@�$Am�<aV��aǭ���ѤV��m=�������01���/���f�V��e����qb��r�s�N�`�ը�������
�����g�n<�FA���^k��G���{2�H7�����:w�n�.蟻�K�g���<����ڔ�O�JhrvR0Y��l02�$�������37���ry$	`Qf
����C)l��
{�/,0�����h�z�&�$͋��ka�Ň��� ���������]ypd`<�� vtf&�K���L�S��U�?#�4�$�g���zΠȫ'�a�Η�ϧsuݱ�k���������L0WAZ����w��2��y��3���̳�e��b�J��E�B���5�J7�F'u���0�Y$���z%���
�kr96.��ᄠ�jc$�ý
.I�tS�a�8��Zc`[o��v�W8FH��F%���ZVo����#�Rx\���l���=r�+��,�o�1����}����0��lg��Tأ;��%�^�����:�g��s�KJ,���:_�1�˗ҺɌPԠ�_��::I��A�����fb7=��UD�)7����\��+�����M�r��8Y7�ŞEm�t�h5#�g�x�����o��h�I��"��C�.]H�͠Q�]F��i���Gm�N��Ձ���~��4k1��:�k���8��oN���09�Ȝ�< e���12�@��Uk�Ef�ʪ�6h�m���O�~��1J���Wб�����F��F^WF�q뉽{]�z�~����T�go��vs����O�W��]���J{�L�i�, ��҄ƛ��z�[u��з���i!�X��7���7�ڥ!o�z
&8-Wv��\�/>��Ȉ9R�Ī~��r'e�\g��Cُ?�8Q��@��KO  8㪩�=��߫�p$�蹳�c�KV1�|�l �!�[�q���!���%#�%�mn����D��&�X����g��P�!2�
�Zg$fg1`����w�{e:�)~6�"|8D�'�,RpV6ӭ'�aV�f� ��0;�>����X,���N�)��qBp��"4�E��θ����!<MD=|�vq�5�(�P�hͤ8�p�����i��A*�����-�e
���O����W���
W���<u�F5�Eq�=/i�ι��!�������A�Ɗ�g���(�jB5D�Lϥ!��~޲8��<���f��������[҆Gt$SK�1�B�TAg0����0NF>	�l4/�T95�v-��A?}�&��цq�W��6�/��;f ��W+	rlS��c�$�I�h�`Q1>��M=���*�	���;�i<�ҕ�4x�`�3� ^y�p�Q�=��s�O��~O����m�7���װ!���Ms9. �_u�&��ǑG�_$;af��F=��m��g^���A���uO�O���$#p��P�c�T�BԦ�p����*es=n�q�v�΢m��Mx�~GN�n0�\Ai?+�L'�׮d�ߔϽű��B�f��Τ�RϿw�n�[cU���Nc���gWӿv��3I��<gfQ���ho_GuI��?����{���2�f��o�{c�Rb��a	���ce��0��j��Ӥߍ,��Y�F���N��Eh�-�� (CS��S`�I@�8"�	Vo���AЛл���z"�'�����x����Yfț��0��킊+h7�n�ge��כ��?�}�W����KZ���<2;#
P����_�3�@l͜�)h;J`����_����ٴ֒�
��|M4���B�pG�T�TTt_?ں��������0��´ <U�� 	�Z�c�Nx����f����gv�����J��S!���{Q��I4�9��=�����t�^G�����_��DAe?�sy^Ŀ�{фfż*ծq�ZD՟ʄ��̰:%�%��q,�p�p>��3I�6��(.~D_��V˂�a��з�IUf�a����`��44o@�(���M�&��A�|�!L`�{q�܇ՈR��FhVM��\d<��qJ����*q�6Sv�.�]�/g��A���벖@ �����D�c��gڹY�|�%ZR�r�v�R�l}�G��/�S���3a܂�hʜ��_3��qc/+���{�1�n�H��]�E��BS�/��|�V��<��:h��x�l��='�EG܉�{P_�-�y,�/=Jxo6i۷G�\T��7x��0w�1�]i�[� ������N��`b��2��jb���S���W�ƚ0��k��^~FY�-�|qbe�������bJc6�~��������#070����f ���^~�_�v��U�#j�/��r��u�Tl��z����+ւB�Q�L���	|B�VB�Q���*+����p�s��B�����$5��*6�AU�>i0���CG�ϛ
?&�9����{~��_�wj	�:�S�d~2��m���r�Us ����rձ�$?�9U{o4��R��x��d��c�3�1�vU��%�����9 1����8�j-��z�",�Dx��	/%[�fb��g������3���e���)�ͦ��n���2���nʳԟ�)X1:�יּ�^g���v��A=�}�w��'>0&�V;|kF`�L�Q�0	�i���,���1�ڧe;��0t@B��8y�O�D�z\WQ��?t�Y�3�#��@�	k��q���
7E���4N�{�j������kTW�3+WTD��O��I-A��<��Ѐ-��~a҂��]$����"�'�����Z���wδ% 5���랛-�mQ�R+���k�gÕ�\��h���oM�{	���لa؄���/�[���Bض6�}��|o3�c\I�+C]�^C0�돐�������Xt��RZ��� �����Q�ɀ���\�aͩ�L�d�ͥ��Y�&a�-ZX#=7*"X�&�S�L5�];���ˊ9�����a�ݖ�l�`�W�Nt��5��N�[c�UO\kI]���=V5�+]�8��{�h�s(��Q�!3�cɒj)Ҕѕ�����G�2k��L�=TO����̏X���G}[�}����g�g��|\Z L���[�Q��ʇ�� 	�����q�$����kə��\�U� I��a̟nzYۨC��	KЇz����[�drMGox�&j� ��zQ���d�%�D\#M�kZ� 0�1Ҋ5�'���uoԁ�3(�#��5��T�`UbE�4f��w�R�x��i��en�����h���sOl�حL���,�*��9��*�z``�D�˳��|$)�8q}���h�uw�#t�������UR�!.R���#�v1!]F�u��EVZ��DѸ:Eݙ	L�>��P- ����Q����s����NG�j���f�ƀ�֏��6}�@77��� �Ta|�ǥ��n�U�2)!w�"����������vT�s�Wv��$��^��$�Мw���Z�Gh�(�0�#��L@bx*#8Ӟvq����ߒP\C�a��2�n��@g���q�8�w�i����::��"�4��}֜�F�u��+���u� ����-���kK�;�	N^e���8~�!af���!�^����7�r%8�nqm�ݘ�8��V�fH)�8��u�jO��c���+4&h .)'�M�q��K�ѿ��;;���#}����������i��Pn�m���m�<�n�5`����I3��e5�A�w��Ʉ�8���b�9���b�U,{�i��$�T�� ��$�U/h�	���O�tep�T����W�/���OM�K��rF9��>�����.����>m�����ag��O��84�����^����Ɲ�̈́nf5B.f^e�귣�X[L9rv��[aT�9�����똚 �������9�տ�(�mp^�������w"��m�
�>t���`�O�N{�i���7�	#�.؝��0`}��%�� �I%�P���p3EbN��h@@�z�W�;n��@&�{y�!8&%2t�hoh���e�м�����7���-��"���6�4�� �q���/@%��sWfȣb�x����K��|������cv��}�Ӏ���v�Vc�}4⠇�@W�Z�\��_5���K�ֲ^�_1J�<��u~Ӻy�e��Kߩ��$�k���6������vv�a��P1�����f�A]��^HD ]l
ʶ�1L��9�hɎ�]��x(�e���M�`	ک��K�r�Gҭ�iɄ���,~ij��D����U����]��L��հ�1ԓ���.vGTG�'�2���S��6�ʾH�":������5U�Q�U8����i�%zA�"q���m�@�7�H�XJ�2|�}�nu� q��������ظ�g��n?��T#&�@܂i|kR75oQAq?TL��~��l-�D�mÐ7�����Wu���?K���Չ-͢�m�<��@A�j�7����F�a�>�+���,<4�2�����p���k<�E�D�?�9�f�R�c}�-7��@6W����0@Z %�� ���_+��<�{4#ˉ��T;!����ZNh��������tꟷ9����Ѯ&Cn���9M�&�\J��vϏʀu�
*���4s���&Qv��*� �Ҝ�7[ĕ	yx�z�d�
k5�軟�H�z�gq�9�i���azñۀlp�-��>gz���ö_D�ZAt��$k�U`�O�zA��*�V��T�G��n\�j�ȱ��V�(US��G슅j+WhN.��8�Jv�-c�5U�^fZؽJ �R]��+BIW�֢֡A֒6�r���݀	��Qzx�Fϖ}󥛛X���!hƼr��u約>GcNXǗ���n*<%��Y��f^o���L	���1��0�¼U�B�w���$V-�������5��������q�
u٦��O���)w�ɰ��jw�Ճ��G?�(s���V�j�B��NɁQ�:ƴ����g���W������"�\ �ȧV�8]�b��.��b ��d��#g��Tk@8,�G4�00�?�;��D�ǰS�?!��� �
���J��OO�'
/hQ�)���cdZ����х��Q��@+,!��n��\}hx��(KjQp���jC��;�w�f�G&Bu�2B�GasO�@�8 �xbsLا��'�=ҩܾ0߫QF��^�{��B��"�vVJؕ��!�`IV�W	�*]#5V]���L�?Bԟ�@eZe-ZT�af��WC�-�%�Q��ħ /�ex�C�&/�ᱩp�s�N���T��j���J�5�h������7�U�^�ݹé�j$Q��+�^��NMM���7�N�n��t�l�'a�2v� �%�@��e�od��ߊm�&��w3�IVF�,@O��Ɣ����s�!����;M��ɚ��f���^�t�����Q�R��Wh�XX_NX����ʶ�aʵ%�󔦯K �3!7��������������ph�{'�i3uk������7%5�I�g�l��WYz���춑;�x&�l�S��1����v>LYk�0�4��m3UbYY��Su<���N��r��  K��ʿ��Y��
�t���	���x�N�Wcց^�m֖m��f�}'\m�f��ǃ�|���;i�D��ߤV[z{�y��/�n��B!���r���{��� G������gk��Y�x��1�u3�����j�e<!�_r�|=-��*"�q6:>Я
)m��R�AI��:�x����?��'�66���U@�t����[ȝ`�})C�]n�Vy+���Y�Q��y��Ӳ��L��3"z|�&���ə��\P�%6u�ćָ��r�$L���)~L��	>U�,F�r��"��u�I�=�#\w��yaұ�����v�q��խ:����:��7����$7�)mu����؁�%��#~�'�A���-��=O ��fj�����?)����K�pz��]%VΦž���f0E:�6�q�+��B)H�`���?j�5�O�)���E���q�x��h	�:®Kh��a9���Ϧ�P���{l���5����\�r�����x0F��LBL�X髸<�-��ɟ�����h ?�%0� ����9B�?�JP�ln0���~7k���ݬ�a�je�:
�f�j�rڦ9����Q�~��)�_+�0�g�݇�X��rϛ0��Qm���#Zg]m�kES�(�<�	�0����Sp����5[��R�2��4��"_mջ�R�(��
��(�ݢe�v���W췭���*k���+���S�=�v(�dȠ�a��$�f!ճ	�ۛ�8Dr�J�1���K�̳<uG���ŀ��OYf�TLI�x�)���i�'�Z;KC���_6�jC$��-�y$������(k JH
�@n�HKc��>ʪ e<�8)��~��Vg��˩ϏEc%� :�h�3�Ҩ��ArB�!_�����3-ӟ�_���2ȵA�}6�����d̊�#��N5rG��/�Ք ��eO��-T I=�k9�/�6��S=.���pn�m���ȽJʺ�:)�P������mf��޾8�����~F�T1��D�eP���5���@�"�s5&��Q��Q#E%aĄi�Ux�_�#�G���|e�v(�9`���L������`q�(>�B�W����sX�Y෩�"8yU᤟�$M���$5e���
;��)/쵾���A#�4wq@U�{�^C��E���<�o�al�<���r} U
�^=��p�@�tS��H�k������+��W�lt]kwb���M�B�������H+�#���T(b-A�)����� V�x�A�T�r9��9P2�FLw�粪&J�����XX'44}h�}�y�|���sDU�z	�K���<��f�(jYy�{0$�F,�+�bq*�{�z�N�man���]�.!�|��?߁�:��� ��Kc��}�A�7QU6�	�z�����0��΢���}�:�쳕Md�ı�Ǒ����5���X2����&4���
ّ;���9 �'z��wtk�$̖(\�g�)�%Q]���?��H��i'l�ZR|��؆�1oh�wz�tk}��L�)�6Ê�;��^��>���B��ܩ�Y�$X8A	�v`֟`C�
��؍(7�ᚎ5�Է�n�.u�,�Mń�3�H��|��"{]�����HIZ��88K�MuW��2�x�!�A�8q��3�R��+�e�?�.M��262u�/�P��������,k��<�OV�K��D=i`�Bͳ��j2&�����Z��YFQR"����f"ذ�vY�7xF	_�>�� ����@)���O-��n<-K+>���G���K���< 0u1	I�k
�w��ϫ���q��w�ot|v��A��~�qʈ	�<���֘����"u�'�חj�!㟸CI٪��Vz�BL5`����f�\�F����۶S�e�v���@pV�,��M��|��	�J5]��'���ss���c�W9~�B�ES]H�H�^N�����W�Y������T�}¦e����R��x�����RY��#2
�eJ,�*��Ю���l�U�5T��4����g����-*�Y�{l�X�Bӽ���%���yS�����?2Un�!�0
�|�i��e�C���5��NΛ����GE�;z惪W6:B3�Ƭ����W��i��(��7��I+�aSZ4��n��lA��h
$�*@�i2"<s}�l)�h8r�į�f�D�ˢRYwvǃ1Wf�M�G >������v���7~�a	���
M��'{&꾓�?�'V?_�5���G�S��V�Zʸb}D���"D���e���D�D)��?'�L�,��c �vw3����Q���-Gմې�Oa�3��'md3'���e��|���n�����%��x���p�ŉ:����&bՅ�~���a�ԓ
�,�\T�$:����>�n��	=s��~��0��e���a3B�}�L 7�;$Dӵ;�Pw�I Qgmx����W���P3�Oz�1|���6!k�&��ض��E�k&fOXi�j`�h�Gm~kir������'<�ps����������N��B�SX42-����*�o,70p]�=���-(�������G��)�X�S_[o��H��0|�W���x�Anҿ�ߠ�+�>�d,�TcF�+��x�wNh�m�a�0��Z�T��+�\w{	�7h�X\���se�����Mf�H��j���C*:�gV��k(��VRB��*�>\���ɹXO�Bő��\ �ZD���H~/5ԹAD�Ȋ�(vx��#����m%D�%T	�r�(�2�>'n0�M��K���O�w^^���ZNM��+,�6x"�k\A�������ayW^Bi����WP|��L�� 8亄G�'�
	t���f-�#H�A���Y�_&	I�5���%�!�z8���Rq����T@�t�� \�9z�)G�/�Jab/��A��	���2�]�Y0o�c�k���PY峏�B�4&>ؚ��Q����0�1Wi`��3�!��S�U!�Mc��O��{laYոh@�3zO��麡
�U�]�^�{n�	»@�7L	Y�`���E�'�v��#�\m�`�0K�� }Y }��"	U 'A��gk��� �1��R���l�~� �߄�������}Db{w����	+g�NK�wޘ?\^�� ۵��l�vq���+��=��F<WZX����^ON{���Gt�d,���M����t皠��m<zUK��h׌W������bX��Dl�#�q��3[�Ç���$P�ˡe��*w6;51>�f1��FC��)��� a������`C�%V*�%S>O�T�=sjz��=<��*Z�%CO�n���	+��0!�}N&g�d�_��X%�4;�m���*K�O{x��$��O�!_g��`f~5���W���I&<>
O6<^���!���d�J}tM2��ӻV�Wj�w-Y��b"�qߣ�~o#���Yd����>����M�AJ�)a\pre���"5�rz2a�V+x��8s`��mv�\��O�Gw���p�O#�Q�A-�m���>1�g�i�/W��s�0j*�h���%K������'��K���-0K�<�|�v�,�����2t�T9����9^IF֒��y��=y�|����0���vꘒ�m��Dnt%�(���[mX���_F�N��*� SG��26ļ���k�?��J��d���9>��!D��"�t	P��ظ��`�C��m����Pf��Z���.!�o�_���r����ʇ2Z�޲D�돎JZZݜ��KWs!�1����i�t/H�12Ew�-{��!�.�"�o�����q�t�8?�sZ�lZ�W���#<[�T�������Y�e�6��(벀��U���x����wP0��*�+�EEw5��(*Ο����sOz1N�O��2�����@/NR��$��W� V���b�Y%��$����Q��>J��3��(+��Y��ゕ��͊�L^X �Z�M� ���.gr�Џ#h�V��V�Ou`h9$)s��Vڌ�6���&�<���W�W��zs<Q<zL��Q��r�aIH�mFE�_"�.���P�[�pw���p4�z)�4;�bi�g�r���I+7|����yܣ�/9F�����T�o`��lWü�L�x��35Z�Syg=��p2�]��kw��#��)�&:�ʢZJ����x�)�i��z��G<�����E2��,�g�f���yŁl���Q�h^�J�>���-F:�?�n�39��E����6c�������S^)��g���ïq�K���uyK�Ղ�2�XV����V�):������M8+N���ә�4s�׬JSbI�"}{]}j�t�!!=^�i��B��z1��Ms_�����Z��[�+4�<bM`+�_�llF����ʐ\�,�Ν�>�dM5{4 �v~cN8鴆��bș� :9�D��/�蜱2	����H&0��ؿl��r ͘)��	�)�8a"��~��I�)	hX�o���N3F�H9��%��xD�/�M?lR<��i/vmC�vT���R&�$_��Y*�~����S���x�1��T���e�aU�t��N>�Z��:����x��|j/A>��-SS9�W2�X� K��*ٙ�� ��FrA����&��� �k��[�x�` '�o��;��6B�]�ma���e����
��R`�=:�w����9>U�HB��O�x�F]<�����5�22��Bp@Dk��{X�.�ei��u8��w����@|���vq������ڕ2���.�WU�(���E�u?8���7m=�\Qy�&�>O��C���!�ٮ�^��+f������U����]�7iPojZ��ӽ�Lt�;��)[ď���%#x�҇����W2�3[~�G��L�c���7�u=�����^���#����dn��y���ed���B�D�U� ��
�����٧����1-<Q@G@��=v�T��
?a�!�7����|���)P��W�	[&��ySۡ�w/9ѵR薋z�H�]yF�ۢ#l$�e2���J��w����OSD���z�zmh	J��s�>�.�{V��	�oc�M�wi�i}r��M��qJ�kƂ:"�1Z��՜u����-��ʆ~�8����"�ǑXD=YX�?mȔ\�w|������e[�b�zڃ^	|���$�'����q�F��D�uy�Ѹ."���`~@�/z�7{�C.���eX���;P.YX�"{n����LS�nj��v�hi�|b���K�D��(u��pj��W�G���x!û�lM�r�TX�*�TZ��{ P<�H-�`nQ4�B0_ԉu���%����VcfN��VW����o�V���W3`��F��]�̺�xmI)�����}�QcüR����4˜�w��el��W@��1����콕�
)��Y_$��sPٔ��7�\�!�۔�$��i.#��M
�����Ԧ<dA���}�N�=j��x�Iݷ5#���d�ڽ"�����foJ�g� ~��#��6�*�HËx���P�{E؞��4��O�Z�E��z�H�0���,

|*,W���9/9��-/�5.���Ta�.3�I2��U���U�W����'�Ka�V���%����_ɪDa���+�e���\�X������f�YR�c�l�-��0����Qn7U���0�w��vK�.{���$���@���c����@s��1�����,b���!��eN���b�9*�kE���2:�ZI3��{H��ʑ'��%���x��d<�Go��o{e��fɡA{e��ܓ��
�s �G*��;+��?�ɇ_;��ߒp�,��z��ס�[�M9l���Z�Sj�olQ����f �R�!Ϩ$=�g���?�a�; ��;}��*L�������n��u�M��K��,]����[��]�;5?b/��MG����Q�lX�o #�	����N�����Ra,�`r�`�g8��̙�"�o/��o?��J���vASu��>�R�oO���![�7����w��3�Z��~��$z��j�w����}w�`����'�K�4���.jpg�h�tا�C@mZ�$B4�'��5���_���S��r�����ܩ--����*��� !%�Y�Ǫ��GS�'=�)���E�`fZ���ӓ�!M�q*��*]#�M�*���˗x�`ۑ�RV0j�s����z��ڐ�?A� 2p}�;M�2��܏�/�)J�5�K�:��
�5�r�"����G���=l��f�s��t��j$U�la���7�����1����j}g��;̕���y���#y���׀1�'[,u�s��P77��L^P�T&m�B�č9q��ê<��ߥ'�d�Jw�2!�I&{$�9W�!1�j�^;����x-����g�Z�x{�Mƌ� � �~n�k��xѻ�����/��j	����d;��� �W�3�(�Iöx<�Vſ��s�[7-+���˸���oq��\�Y�o��6��:�r �ߐ�K��ʱb+���cX��W{��
��1�<Dҙ{o\{�%0���'��%�J�=|lW,�q�v�/ҳ�V̰x�E��ZO$VL�#i�U'D{s�,+f�(�&����[k��� PȞ*��%哖g���s��릸f>�ZGOs�Ԏ�<�+����s���n99r;c�CxTЋf+��LZb��'E�c�h�Ur�xY�BP�R��h���@uh��ȶ��.��h�+JŐ �hW~l���H��b�r�A���(?
�l�(&)OS~ɖ�����g� ^��j�0�aE����d��K���Ly�� Ζ�
|m�f߫*	P�@�.����<�������&����WIJpf؏c�"�<�R�i�V�!� #<�������Ҽ�f�@V�%��rs�����t�M��[L<��[�,(ݚ:�r�ù�gr��|rb�>oIJ�kڕ.�٣S�1�w��� ���+��i�Om�q��@�UcO������;�,^UY����46����K���wjLσb�H�o���HUet
U�{�rp�O\�wU7uJψeq��F���� ?`�6k<#l��������w��$��0��0j�^?�T��hl�.� �|N�F D��o,EQ2�]��Y-}ekZf���d��Y������!�-�DA=5�o�Q��2�JZ�?���9����I�0�M�\'�l,cd��h�A���{�յ�x�+~����Ѷ�M��9:���NK:��n��ʯ�_m�dC�-ma��UH;mW�����W5W��λ#f��8���L�%�U�H�������D�W�n��wD�CS:�����R�V�אy=��A�|7��6I�"����6�0�dʺ(e�b&�#�Pjŕ]"��nۤ�z�O�+�B����4�kޫU��_�
����+��.� ��3��(��j�h*ow�,oR�oOۢ>��n=R	ܖ-�܃[����4i��~H3��(�m�C��b䬮k�݊h�[�gAn�C�T�����N��u�4�9	�vjW�'N����<vC �̓s�9y���Ӯ��@�a�Y��U.D�hjNN��������82��N�)�|���8pp�P#r-�u�o�"%t� F5k�����b�M
�����Eʻ���ڎ�_갤��@��\Yg�<q��:潉�"�`s�Ǡ�^WnӋ�el$wc�Mt����H�;��=.O�9-�bΚ{��J~H_�%P	n�Hhx@&�?{e��!�0��ի9�w��Q�P%X��*�D?4��ʞ�10���p[�BQgIJ�i�J��;�XZY�FZLt�r��1��H�����cl�X|L�h�Wh>$�d[���okQ�{��ܓ]�|�0�*-�9�: \��&���̨���9�u�([a4�ڇ���fR=AW{М�E����n������e�>�}i���m��ߴ�Ts�L�Бp׳�mA�y����/���98�X�R�ԇ)�un���t�h��B^R<��6g��>0$�̂�-��]��sy 6�p��02O;ջ���Z.�u�e�-S���cw�; �ώR�-�A�1P�6DB~y>R���*>S!o�ʈW��|IT6�8��)ل�������ܛ2/�a2��j[	!.���+׊v�iZ���Y�k�:�:��q����= ����8��6Zu���ι�p\o��_�͠j�B��g����y</h�Gצ�%@ˠVn��# �1���ԇ�G�Q�nu �1����@+o����Ӝ���ɸ���)���V�?oKu#k^�����.9Q�JB�ʭP{h�g&���p:���t�sν��ڟ>�q��
G�vo�֍��D�t�:�;�h'7��*�?Yڕ���V3�/�ǟJ��3�5m��^ ������R�p�0�0������"��ka&W���������mR�+m|�]"��&�d�v(j��0(9�89�z�t����Ge<sQ>���q�k<'��u>;��>���H4u	����vI���T�[O�v)����Y��u�C���[�{Js�������@]��Ŀ.@G|�C�Q����"�z�cE>i`��<N���\���*����i}O1$C��h`�.����n����@j�;�9�T'�Q)N�;�e5].��V%
P�Y��`U�Ax��c�����gz�/���o��� �*#w96�ƗX!*��^����Gn.�j�*��u��g�B�|W�8���Gn.q��FU	>���53��}5�̩����l�"��L��(�io�"�ג��>�n�G��j>K4���5������u��ZQ��ށP��be�|~����q>i}0�(e@�,��&y����mc�XQ��_�:Z������Q%st�����2ɹ%��f���j�]�&��a���>Q�����4^B����W<T��G\|��,������>�1�H��x�5�l���j8����X�A�1��I�L:-">��d�)DwLn<��S���L#��6�~�q^!����k�n��%�}���*���m+w�Ui�Ċu�_�I��",t^D�v��@��Գ��M�{���{E�@"�%Ķ�iLO2�l@!F�KS�>�zj��vpCdw-�"�י9����@F/���~��8ϝ��y�{�cy�g��5�	mQRj[GU��1yE�߈^��¨�O"YA�&E��
���ε�Bb�J�)���`i����_$߃���A�T����t"�m�*}3�"��=HtrD�z++�3K�43��2���Cl�!@����c�����rȥ�_.
d�CI��W�>o�i��p}<�qV5��/�V2�.�B�,���*��>��+bo�w�#���K��/ $y1�D�1�τ�:6N������H��9s�򃌶}��`�8��,�zn�n�8/Y�:���,������\�E%X�{�@"�5d�.�i.4�������z�aj�ɦ����^�^���!Ϻ��b������i����uX_��h"�M�X!�9/xDp�!�ca6�׻h{V/�I��Vy=��l��m�$c�;!��l��9q�l}L��pDq��g��3�5O��T9<��6Xp��3[�����З.��R��G1�oz�tRʮhw6�pK����x�nk�GNM�!��?�)Ů��D�a'��uޛ��jIN����	�x��+����	�
������/��|j��˨O�w
�J����$�����|A8�Y�3(�T�����V9#�;Hrruԁ^��܎$��TE�Fl��f�%��`�D,w�sG�	bp)KЃ~�a+��G����w1$c:|�ow�������&M ��O8=�>߷ڒxX��� ����|����k*�B�����nF���vT˞��>�*v�}Í�A��#uR���k9&�����/�<H��N�(I���}�T:�,g���!���x�"հƅ^�ϜB�ҧV"�U�Ln๥s8"i�����4�Ĩ�n��#�1/������+o�J%���F���C#��F��H%��>`���-3���7����c�M��2ģؘ��b�$ ��|lt�*�G��c�og�*h�Je3=�F���׏C&���C4�������#�CZ{�"UM1�<3����%��єo�t�nƜU�<�*E?��	&�/ٿ��V�z��qZ�Q�y*|WI�G�81*���&��X^����T��J�*~d���O]�d�"��3�~1���*��ڮc$�3��� �T�1�}ڛ1��=*>�|l���*���ބ)vͯ"��X��'t@5EM1w*�� w���A��j�@���@��7c�!r�N/u�L�N��R�n=��#A�2����q}�� ocȂ��=J����KpVaQ�%�zo���U#��אNoF�]���5"H��I�7L:Jym�
�`�G��v��+�"nE�V=v��+c$a��󟳈�(� ��1]W���W�D��� ��>m
��@��4���#3���w�?��˼ �����y�'w)s>���G%Xfv�H��z���l����R��%����m(�6E��zoJo�TWh�F>n����y�JkꇠC�DR\�T-,��&ӭ���i���ܺ�\��x�i�9�D��� ��;B�kJ�5�E�L2X�v�C��0l���vExx��HXٍ�r@|s6�v��E��1�ef�_4�,��?���݊�C��U�D�;�Ż6���lU�rڣ?���Q (̶,Ƨ�0���;	��T?��y[�7~�Y��B5
�N�L~abl���skv�T	�}!���Db>|���j#� |������'��"�ӫ�F$��:��+�Y^-��IFF2�|�����#� �O�Xf��z��&�Ȋ�ƾ�NW�'+�r-g�֚�������yi:�kH��|�7]�B�|�p���l����m�WY�4�1ɘ��t5�0 �Ӵ����>�Ǔ���Ymf���w�X�`ݰ�͙���b�����@b�5��^SH�4Aн�V���[ʳ���Xː��S�j5&� I<M��#*�]�U�*�ã؛*�*8��@�8@e��<s0��df��69bu�����P���jW�U_�B�c���(f~��	�ޏʝ�K��!}��+v�\�	Y�2�ł�)�A�c�T�L��l�U��` ���E�W��e�|�к@�w�>hr�w�q�憂���'��R��LSG�U���~P�;�v�]�Z�O�@���܅� ���5�|�ҦF���л�2�o$����a����]��]:zX�S%90@{Hѫ� ����@�I?���#��p���k,pPb�� �Ƞ��@��z�~\I\`��{��&< )B4Nm�	��D\�^S��N�;�c��� B9�nD���#̎R*<�7r��;�e�g�
�CFn��v�	p�����d���O<=;��3�`�V�j߭�=�oe[wF �޷M����F �`��|���uI��UL&u��\U֊���f��\�� �}�w��<|��{�]�Wh���iJQCNy���lGa���,��T�T�FY@�΃�������U�����X+���}��SA�V���t:С��U�0��U�4Ю�{�^�`���To;GԛC�]ZY��Y	��UJ�f��1f9��H:*�r3db��cѫr&́�rU-�K���|6�iԅ���K���o+�Y�b��"��/&�gE^O
)�=�q�-�妣��������{H���@�.]!N�h��9?p?s{�U�z�^K�s5t��W��߿5_a�
f�M�#��/�d�"lѯ��L:�`}�:�Q����đy���#f2�����6f�S�'ak��~�u��;��zǹ# �dJ<x4����!�m��Z�4��e���U~0t'��Th5���G��4^̌����l�1���{��\v���'�}���2�/Dx䲉9h}
��ՉZ޷�$lV�9�(����|��� j��?%(�?�S!�v�D���.&���m�)&!�AJ�,�UEg���cdw��.��i�rG��B>#�KT���א�bc�`4�(}��B�HVm�����8�[���5MC����-24G	�yθR�e�\	BG1��:@��l��3�1���b�ZCE�{����zF��ψ���Qi��9�����߭R���-X�:Y�?S���#PC�z/W��z}�e���LHx8��Kk�g}��ȺH�Ӣ�
5#$P&��h*c ��KӒ�φ㱃�qb	���JO2w��"��zi&��F�&�2p��M�� <S3.t�h#���!j�xnz_jěҏ�U�ǑYK����6(k����	�TPYv�ʍlW5��]BˏA��/��=l��GDC��������s���oLj��I`������_��?I|�)}�����v@Tvh��Vw{}n�t�j��&���NׅI�]Vu���o/�F���F�uo�����9 ���>}���"�A��w�n��۱hM�F]L}_�l9��*� ��U�3{�'^*@��x(`zg��'rA�����M?L�����p�5�ǠWI��5�6���\�gh]Pnd�M�;Hi9�l�dq-�N�t���\	A�o��n�)���(.����Z������(Œҩ��SIe�2#/�U�{lrA�Z�A_�|9U����5z{����!��@���uy�IS�9��|�,eG�le�����i���9%�3���U���5)I���`�p��L��K�\���7==1K&˺کf�\��{_����,�
��LX<��if��1�a��N�P�+<Y�z���ϓe����6�P�X����坞z}���_�2�h�q�{ͅz�54���W���7��H����]yb���Zf�"�YI��?���O-�ö��3.h����p�q�t�A�$�X2_J�� ��L����j�Z���蛞@�˧��ݱ�ŴHңD��Ŗ���$A�v�"0+��}��G��^�(�p�Ca��Zڒ���8����b��	+\F�H<EZoPY���٣�׸�"E3^���@7�W�b�M5=�Y����y�A�6��i�x|���ރ�Wn��i3�ޗ�$�]w1ָKg@�]�A`�.�奤}9߄�!�U��]V�t$�	n�[�a7F�	7Z�>��=��M,�O���0�� :\��_�
k�p[��b8�=��#��*�';�x���nb�l�s��zҜ��+��T�������$ ��S��ۢN�;�h�$���J��3�g�*���#nD���4�\u-�2xW����7�tv�� :m����ߍ*#�"	;la��;|�*�xg�bz2�'���~�LȤf�ɥlZĲ�n[��L3;ɨ��U�Ȑ�Q�� �ty�^U߻�,�
�|������	[�'3ψ����V_�A���qӂ �DLA�,��
��[l�;i����+�fT��H�H�'��vg t3^���ߒ���ɳd���ޝ�Ή��+�8)D�+�=�(�f�uJ�r)n�������$�TY�lٓm4d5�/I�������æ���<�Z_�]��SĖ�{��� B���j��p����;gg�^�b���!<�0�G���f��I<@�@���r���t03q���{��}v>��(k��ճ��N�L�O�
m�9�0C/���Y�#� �n鿿��.��L��j�!-��fu_�!�f�t��}��� �{#����\^9�ƛ���}����L������������X�޵���`���>/�r����!����QL�W��{4m���D�abrG�m(pj��C�`Aj\���8(J��y���U}"dQ��?WC]Ǟ{Xk�PA�����9y�ר�{�N��G��ƾ^$Kv��3:���w?����0�4�dϞ����`�*3�ގ�2B��&-�*�ӑ2D��f@�٩��)���2h#H�ES0V�5}�lC����Q�9�@q�L������=�r�>i�S�)�A�X,����=�J�!9b���\���~��7���}�y��t]YR]���i��6�����<̬yZ�����M<��,��mGF5��qs����"�h��d`u]�ס`�v�*{1)�Y�3$����L�{�<_=$ Q\w�ﴣ��?�k�W�]�K�T��h4\��s�&l�� ��/�8��Z���� 㶆?��f�υ���0r��:uDS�z�W�d_,�Q5�F��f@ޑ����I��'��d�½W�?p�kŅ-�}�N2�bU��zc��N���؇��:�К�q|6(KQ��NY|5�!u���ar�#	ǲ�L=]�`�O�����N"���ՙ��<����&��&j䧺��;\�ͅ��︒�����5#7��O8���+#z��X��c����T��=�~�㟈��aM����x2�Ud�跎�FE���7&]\���4�7ZF�7�|��$qi|�6�7�_Ij���Y���j�Lr*�����u�n¦��X�4�I0�F�M��5i��~����R���^ѕ��*U&�;����Q��YJ�����Av��Y	~�M"��Hц�6F�D�a�c!f�2�U�f��D�/�28ODj��s��T&	WE���N��޸�y˙N�6�tئ3{�$&	h/�N��͒P�����Ȁ���9�pp��]Xoo�
�c���3��m�2 �lD���oD	�i�`F���������v(H�|}x�TK�`���qӉ)��I�֏�J�Ծ-0���Yra���k�M�ϳ{�*�9�>����Ǩ���\�<|����;��n�~��W��+�
��6�2��1�o�)��8���'Y%
�Ԃ�P����Ƞf3ъ�u�i7ШE|r�3\�v�ws�?�e�H`��{��ֻ=�_��pt�͆=Ůq��/-�	d�E��x\A1����Py�9ΧRV�2�X�h5~����C�0࿫���h�
����?�2i����fkc�n�}>S�T�-��X�"�y�?r���5��+�lA+k��A�5�Z�P'Y9�I�����/�p�v�v��%��%�TW#D���$>7yT�J	�3��0�Cl�<�i$	���l�[�����a��_���K�6CB+�^�������� �����_Yy8�R�Q��|yc�����2_Z�M�)�ʰ��i��[�ʍ�jvA�֫�	�p�9k��ʂ�̈!�B���=S\E�Xϊ��yx��[�yX^�\ YWU˵�u-1}î,�`�]�������*����,謃V��kW��
5��%|���a`�������r�={��3�U�R=�;ϰ���&5i<�-#��	zR�����w^2;��"��~��[![�9!i��(Ip�����!��׋�"�^y�䤙s�?��E,��x5/����Ze�]wf�*����U�T[�j�r�%�P�-��`��Jx�Cn����kW5��!�UG,���Q��Gb4�z�`�-�4�������U��菎߼N:2`qؙ�q�j'��MN����\��Y�ă��{T�3,�tK��YQe�#>Q�˻���dߡ>\�Ɔތ�����p��`Ҧ�Ġ�r!*Ȳ�#B��ܩI��Z���Y��^���Pz���W^P�p��J(V�]I�z.k�%���ٷZ�60ul>�}����u'Tʄa�����⟍M�v���4	O,t��4��,�^�4Je�-\4ke���5��1���ޅv�byi����:�B�����(��S��ە �W�|o����Ƌ����%��X�!�a�rv�=Bz%��SZ�>��;ۖ�0P�����C.���Qo�%�W�;��̴n��9���d�a� �A(Н@�y<1֗�z)ށ��5jE|A8r��B�ڦ��?�+Q��Y�u��~�����{�.
���R�O{�����~SFя��1�C��ut��3\����Wz�9F�6����� ӥ�QX�y�.udLX)����W���g��r��6~2�;��-T�*�|���FG�Y�W]�����3�"��%C���B�3r�D�
��ݪ�����8;��r��w�,�e���"U��;��l���O��-����@�c)p�>�U����}���Y�50�!�IjE:�m2���'5o��#����,�3~n���N c��c�N�O~2��ɂ^�-�ҥuv�F��0'b���j˦�����it4�8dC�I8�ʙ�Ҹ��t�L����g�ߦD)�r�\�q�Q�[d&�+�H��:��J��PMȨ���ti��6�

r�-�U���ؓ�×�������Le���$oJ��Y���X�Gژu����w�U0f�e�c���'X!i�z���5{��˴×�Q�i���~�(�Y@���lc���͌qQjy��\фxPQ�,N#������u���"<� וk�\ˠl�g]��5'��]�*If�T��hk0M�;{���&�u6�����TЦ��A�L_+е舴�\�&8Jb`�leu+#��Ȏ7���p�4����[��`9�'l�xɴ��c8觗٬�g�����6�L�e|e8w���n{*��S=�p�"x�La�[_�����4�g���͟����#9}
��
�Ț>�R����
C�L��������.mz��N`������T��=��L���P�'f�zo����a2H���i,VI��d	5V�#�fbS��QUD����o�4>CYy��>z��6cO���-�mbD-	ɕ�mtx�W��c�{Uĺ��*z����u@n5����K)¥H�3��)3�T>^̮�dTr��@���z<�,	nB瘓�X�����๽�Ӿ���\"�<���r+}��%u#!ƥ3��ↂ��j�]�˒DU�z���&��u�:�W�㗜A)cn�M]t4VԈR�Ӑ��F�B0CNGӆİ����O�\����v\��e�n;�ԟ�������LW�����=��{$)d� �j7Qg[���{�cFm'�e���z��aS��¶9�\��ϩ��R���秡�K��gn��^"±1۩���DP��M��1>/�t

�嫻'�7[l���!�e���@��*-�.nA�]+����:�c/�Ҩ'a�a���h,E��FUlW���{�j>8�ɠ�BQ*�
ϟ?	��3�D��xv_����IP�QL�s��E&<���_:��fg��;�z�	l]�5ր �	i�"�"k��S��t��h����2�K�*��[;���*l�������6i�-�3�9U
�rx���5�DiL��Y�9�G}���b� 0���=��Xn��.�k�PL#./��d�Ӿ��+���g!�Ĕ�o��e�i�A�[P�� �-?n�.��=m�c�ж�%�<bWҾ�[��M�M�g�M|�����9\���ʹxr���S@t����y���\=��]���H�Aj80���k���c��d��#�4\*?�fH��5��Dgy�0�q���[<��z�9�|�}.�M�ΑӪ�/�"�nVrP)�/*#�i����Q�l��g\אK�9'$�`��8����t��ς�{1F!�֗�V'-�$�6e��Fk�����#��]0�i��G�B�X$ů����*j?Q�-P���X�/�ᙖ��
V��xvl��W�G��aGoҶ����
�mԪK
`M�K�E����{�}���UӪ0��K�O�ДЀ�N~�����V��	���j0*8���]�1�ҢγBl�:r��J����N1d��LmV�*<+o�yc���b�Vto�s��D�@����нZ����S�_cЇ6/�7sB>���r���O�G؍�fNl:H�bD/e�8�ϩr�wi� +ho��n��kҪ�I�U�f�[����Z���˾���=��=G��jjv�M�Z%$�X9�^>��虹�*dF]v��}�,�b�+ڞ��
�<�?R�1�D��Χ��T�ɒ:X-V�9��2��x9!S�k��{T�n;@ó\��i��"&��#��.�-�D��T[�BP�tif�(쇖e��{ �v�+S��>������^�G<&qһ.�k��7|�nS]X)�a&?�rx����O�/��2���%�?�@�%}� �Œ�uo�!@���~C�)��=MK.�D��Et��G�iH(�R�r7qs� �y�B���u$?����X���@k��ʀ��ۙ���85��E�#���ú����^�a0(�����I�#Uy�W��/��N�����K?�U�����/�� Ƞ��"�'מG�� �b�
�~ȫ7��W�C�����T�����ܛ�bt)r�-{���V������R�(��=�Jy6��hrF�0ɮ�^��J�r6��z�z�z�9����YZmͣ%m{�t���(��!`P��e'�^!�
y�ؘ%dJӾB��ב�z�)���s�'h�FP�Am�1Ӏ��h�� �I 5��!� 0S�Ü���jC��sIS�A���Qb����_�X�p�s�ٵ��F؆�]�U��b��+G����b�:�V�L"�n�%ځ3��S�z�a���P��͝�k\�a�SL�Rh}.l2B[Jqg2�y�_?��.s����a���GA��Nb�V٥X�4U��D�g?59��r��f(�*B�ϗ��%��z� :��ʾ�a�d�b�a����!x	^K4�/�{���2����a�"����C�������5�iPxy6;@�1l>`�e�I��XE�/�܍*�ciՒi����2D-���r�"gV����MB��O��HdL��0�ê<U	��r�W.����U�NߟK*s�p������{_KN�X��_�U�LS�T�M��q�GE!�k��:��|ُ�� �>��Ã�ᷭ��yH���p�4	��F�ӓ�]KS�#�'��ds3t��i&B'�H��KT��n41�8A�?$�\ �2��1�-�pVϚa�p��dǜ��.�תF�\�k�8,�f��@������[Bx���,k��6
�_�A�0ʟ5xZE � �A2UU@�3����+�C_��� Lr���#l�x/����^Vw�)\D̈��B�3�bO��u>X�}�93SRc%�[��"�R��{+��K��U��Sh�]%���J �$ ��d�)�}gNl��\G������x�%�A�s������j���ԩr�»Q�%�]&�}3��x+���L�5����7
��V���&P���U�x��a̘��
���� �:㾟��\�^����V�K��viD��ĢxCL��������_�01Չ�bx +�ݴ_8^е�q��XZ�]T`�h3���V����'��:�B�[O0d~/S��!��,�X��[�ԅ��$]��FF��y���x%����ccQRo͚�>k|������+M��v
7�o�O@��>�uߖ����4\o��F�i�!m�=b�#y�b�b������W�J�c�y>K�1P����?�ˡA =���u_,D=r�K�k	t�ǟs�����cԡ1�<r1�]�tk]u9@��o������uϳ!A��[���xK�9�U1��Z*q:���k ���a��^�(����ss�z6���A�'�,oo���}�$���[�6�`�7����S��"��z�V��W+�2�ި*�wȌf�\�������~�9��;Ѣq���Z�G y�$��U�jY��!ꊮ��!9�5�{�2ʄȫ���T3��KJ���<�,��{�:�$�'4�i��q��55��=�l�:�ߘ��{rB����1ԶZ����sA&�|s�7���=vd�x�'H��뒓�l4F����.A�ȋ:��2��r��b)�dD#UȰ��6�w�C@t���(�nc�TV7��Lp�$:,L_"��gp�"�J�grF��rs� Ǥ�}�S��_*���r?�pq��J�Z!%]�H�f��5Y%m]�ҋ�HIOu�^fv��l��S2YX��#e�(m����`Q�:���bCQ�j�@_(0ݷ ��J�1�	�:k��x���6�^P�?f�[�gE��l*��k�oą��T�֧���A|'h���9GϷ�`)p��)��ҧ�G,��n���K܊/���;_	ZFU3��:lu&�M���\���Gt/��s�/�v�B��KF���.�ۼ��xaJ��ԥ��w+{�O^�G�ɘЅ���z�^�|���(�;��QK8tO�WwK!�ɑH��~��9Q�c+D�i�z2���J��lވ#����3��
��ӫ�0}*Ѐ��OYé��������4굣'�zú\(�&����t	n�Do)T�Z� ���/`�Vdc�z��&r4�*A�WQ�Fޤ!�Ǽ��~��j�U�!n�\��G��X穈��t̷�@�=T!�FG���)�6����Aq�"H��݇����>�>V�Kc�@�����6Y_]���]�ryQ�{z/�#1��OmԮ��'�n�a����,�&�W��/��^�uL=�Hs����B�ߘd�|0\~�	J����4乍}�鹗�
�O�оYq�5�l4id�L󔸨�R��������b����x&�Ӣ��K�舕��%��%�a�0��c� ���֦
��[�]��Gʢ�������ϸG2R���ۊf'OF���[�Bu�t��%.u�b�Q�3���B�(ڪQ#��⅒;*Dy�z,�~���L��i2�``|0��(��,,3i���~S3��_�"	��ϽdB���XT��5�6����֎sT{\Q���T�������Nm�}��b
|�Ea�9���������R9F���\闛Sڋ��#�md4�v��7�<�i��> ��E�J�JQk�wQ�2��I�h��E~���O{���'N�k��(�]0��^�����_�-4Ѱ#d��7�d�ߒ�dP>לb)�B�W�V��=���yR�mv|s��4M��m��Q�H�֝�`.?;�����r=��:�����1���G�Ɏ 5q�ZP���~򱽦"�� X������I�E���'6]��3����bGy6޲���m#l�9�ȵ{e��'�5V��!D�
<O�.��}�~h,����:T0%��R��"�6]#r�*�"�h�%��B��)��l˖n`���
��3#��]A��Cgu N��p`�����^1vX����S����fµp�Op������63#�2W<|냡ס����#s����,����=.bD��el�khF�b#!ӯGy@�$���[5�T��	�e��@܂�y�و���űՂ� Qsj���_d¾��� ��sS=���ѧN3jxf���qyRrg�~���Lt2��$�E[&<5���CĜM����O�x,^U����!����J{����H�j���#����~���=��U˃z�1y-���R�䂣��(O�FܺM=*���P,��N�g�o,5�^9�`~ +�d��i2,�����\S	J��.Kh(�iL�8kb� ��=���)**7b�.�׫� �Z��:)�C��H�|�C�F�Z�k���VL��4��O�P;�Z�`v��@�:�.�**ey���)J=�������n����:����ƺ� a���%I��1�93R��k�[�=AD��Y`�M������1�@:�'d)OZ��ov�����p�ġo�_*��RLV��%
��{�ry�����rE�6����!���(8-5��⽬�:���p�%!Ews� ��OxE�R���d�p�V\pw��`NlvK����r˓�ܙ#�6�+�v��(r�-��0�K���{�ChS�!������$�RF����
gɒ�I,��pU�s�����$�Xt*�$Ck`��Xޙm�$��'�l��4dc�#Ӫ��UC�uJ�B�ob-��vZ�S��c��N����v5�?�`�����<'$4tm�Z��P�'����[tS�X��b&&��@�7`4_���
�85�����]�K@U�������o���_L5��K)��MQml��/7��[�_<��{��@���nՅ9�:#9Ц3��o5Ol�-�R��N--V�А��_��}��C��u�4o���U٤Nҧ.���袇��w�VTSa@�q�|�1�Uߖ���q	�K1�+���k�<@�����թ����4H"s��ގ�Y�z���ByIc��q N��������\I� AF*�_ĢI�M�Wz)�'��oz�y%�i�9�,CqQ��TWZ
�� B)��ё<i�ܔW�~�+�����<y�ւ���&J���=��G:
�b�8���}]�b��,����/Z���v�� ̨צ��Z5��n7FO��M�H�r�����{t��[5���Xz�]�`��+Y�AׁY�����`P��9KΛ=c�l�**���A�i� d!!Ҧ>v�7���cw�i����+��$,/|�cy���u��,,UT�{��^�q�Cb�+5M�X'���Z6A�&Q�}~�����W��[�jI���VDq�2�R iY�_��	����'�kק���G�#Η*��LV/��([���ܿ<j�֗���P/H������^zt�nt�a�\oǟ�x@����]�m�d�N'aSWjqh���4�I�{f_��E4�|��"TRE��"�*GG$��>s{�f�	6��]��Ht<��������+��S�_��Cc'����۞��|��2��]��0Qz�Wd�����u
���t�e:�|s,\m�>��ydcr�awm��y�i��d	c��y���1)an� jY47��w�~�l�%���-+�<yQ~�qUB�T�)O\������X;Y�hk%�����w�{����z��u嚚�����;j�k1��&��$�a(�杒��Q5�)p=8E}��\i�]ڭ˩�������\�����c�W��6O��>Ř>�Q���z�*���l�P�o�`��6�iGѝ�����4	x┗�]�HDWW������� g�@���T�t;�z�3	S6�K�F�L���iw	e����G��u胑@< Y'g�c{�t	�Qs����X�8�+?˟z����1��5��w���g�FniPt���s��z%����{Y�qF�aE6�.e���2�o���=�t%�k��8�ݲ���0�J��Qf�t~�Je���ػ���mZ`�oPQ��Ejr�s����x�P�H҇�p�{@F���2�����d�����kL!�L��lt}��Y�-���z8ItO�+#��1>�M'}��l���*��Bi��"4A�_�A��yL�R��	@+�Fo�v������<R�ħ�PZA��N�G?�;/ ��x�}ޣ#nL�=�b0=��$�g����C�Z캮ɉաD�(|q" `;?8��ވ�3�[4<E�����_�8���컪IV$�������eL�XQ���ida])zP4D~3�$�:������w�ɋ��r���J!G(=�h�F̪�Z��5>����'�(C��	$H��,�A�خ+3[	���A��-jp���u/�'`�6[B��@��m�i��"�e�T02F��~���G�O������{��a WDj9E
.�
�/��;,�L��P���F�2XD�Hy�-v(�Y�	7���]��=
�|R+�}����@LhJL�鸋Rۊ'�!�y?.��cY���ɸ	�D�HF�Q�({�"��1�qOb�����Q�P�]�KM�Xs���%0Ɉ�Ri=	5��7z�
x�Z{Z�'�_,��	�n8��+�\�յ[FOq3����_B'����:�l	���L�I��,��H@E5;�pM0�Gp�
�3,�(k�0AŢq;����UC?
�?\��?�<�ھ�
�J��TH�)��D��au�]�̞?z�,CrВ�(;=��؊��z�E@�趩�B�D>.�Hr�>V%۸�:�`4@�=kl��x	�]_��k`p/7n��=���ҷW��8�P�q������������2W��DՌx�i+���?J�d�d�ǜ���P���+x��q�置�п����O���oHˇd�;�ݎ�H��ٝe����}	&��9�*!���ȊXbZ��j�Nb9Q���w��N�v��He����Q�9\7��+8�Z��@4���WW5�i/o�O�R@[�`����І���&�� 5K����٣o�eA������>)A:2���	�VI��:9Sq�O�p6���1"���61;W!�&���"�V+z�V�ݞ���.)�h��>DP9��\��4V����I	ֱM@�R��eL�Ѯĳy�����l�qywǍy�Jb��&;�~Z2�x��i(�#�[
���Υ`%����"�xM�O}�?�'��Jo�����7�
�WN<HJ��T�����?���ɋ��i�T��Q}�H�\Y��ǯ(ȷ�8݅0��
I�WƂ�5�*ѹ�q�VJ�m^08^�\;����ۑ�.p���	�3� ��L���i�ϔ }
��TH�oDm��򉩱�	KkHk���C�)��������ϸf�b�Fê&{0�[ܼ�Î�`�!��I� ���8=/Gf
�LO
co��w�����"�Syؐ?�Eѓ�ήu���Y�dc�p��)�(��i�>1�<����풻0kQXi{��ߓ��R�نT��V�@����e��%Z~%���;���_^j���j-k*@�ܗ@N����?�ǯC۳\[�r�������s�v�*΀�`�>8|��v�s���)�� E����6ڞ��Z
l?�F_��}�HH�0M+Ҍ��/���;����y�@NU�(ʄ{A�>;A��i�tv��ؓ�dD�|!ǻ~ΊYB�	b�@y�F-ݎvX�v*�U�i]�4�Z"	2ϸi�tS�P-�*�g{���,rº$*0^ӂ+�Y8���@�2�$յ�\��n�Ef>�b�f�:p-0wۥ2>�p.���cd�M��^.���!�O��l���P%��6
�+l�/)���g�-�D�j�Y�]�m'���޳_���zV�f׾G����ᯚ˙A8W3�z�=���|u��������l�c��ؚ�H�E�1X����ٖ�/3�=�f��K7}�%�|΢�� �jZ���1Ԭ�9	�Mv�DX*�@-<�E���ch�E��Ѐ6,��C?5��z�4Z�M��<@��J�NU��t��TIHmo���C��N��^-o� �o�ˮ�B��'+�~ ʪJc���(�j���[�GU��ֺ�f��9"��*\��M�=�,蓏�6�W�~�2�T����+T.�889W	�\9:�?�@-#b�e���1c���X�W�����N��-�|k���Șs[V�{%�á�2c8��Z���6(�q(�QA��	��U}�v�'s!}?�[��ݎ�')�GCvh��vpZ�zt�*�@���uA�,�S�~�I2��۬�9C�`#ZR6bA�-�.ᪿ6GN ��Ӄ
��7����h�s��H���g��Q�����ſl����?��B�w�MS��Z�!U�}H��a��̣A��n3�](�ȁD�>����b�Z,š�G�L �k���ʞl��;�1���Q�]�A����
ۧ�L����Ţ�VU8�w	����|Ď謁qT� ������i��tv�<2��)7��J`*��^��s�f�"��c��{>�"�ͼ��u��a,,p�@�ɛ0�EG����.33{��@$F�){\���2Qtٽ��/���(,a���X��"r1bZR��5��5�jT��aбG�膀��}��s>	�Aw��L\n���a7J�E��Ւ-��0���U�<��QeLo��y�ړ���.��zf$x�ȓ�N��:�޿fn'�զ��(a�{��!����{��9��j�r{�g;P���D����0��	.eh���,�*��}� ��/'�ԱN߉Kk����#	�z9xc?��)�UP��̆S���̣��k�R�l�CѨ�!��J&$�H�O&"��n�?z@O��-��I�>gIN���3�h�/�����,>~�}�:4�_��g�E�I��O N2���	�/�Mu\�+�!���~����5J�]� �5LJ���煛��2���0{��YV�yYV���0'�~����e?wQ<ޢ�)2?�%����\��dY_��R�U �&�uE��H�\N~�
;"KNZ�X�	!V���L{��r�d���3{��Q<e^�^c8��)70Ig�v��DT t�.1���(7����[�����D��l�����/���e1r��jzq~A��9j	���5�m#*2�$l*<Z�ܝ
q�3�m��T7��]�/="�L�|�9�c�u��&i�s�&���>{�*�	(V�$��o5>�\�,�ڰ'��V����0D�}W����?%��Dì.�3��{3[:��RW�N	8h���I��U���牒1(�i:b�Gq��-�S̍<2����T,���%�R��.b���X�Fb�l&9�U=H��s}OB>3h'��J5�F�ciL�
0s���d�}��-�2���L�O9�u^%<i��X���/;�/͗��w5�
1����{z�4�aq6Z�[U@I�# ��wk�C���54�-�!r�v5e9�ʬ��z�~��>4�_բ9Z�s�9fըP-c=�ĭ�gnԳ�|�$�n�,�����)����O5q��+.�&?eZ����<˔��+�|���'p�=ʂ�֑��#��(�g�8k���R;�l��2�����?c���0��Z4#P�lqZ�[��h����M�����+��C��«�z��F)�}� �r��"��h,�1��0��+� �7�v��V�/��V��5SE��O~�WC1�.U�ɚՕO㫵ݞ�3��N�/ >7��hJ�@e���%�?�g�F9>�b��]$w�@J%�=�Jn��>.�O+׈hM�ѥ�^�ebA)M��⭘W�}�1�{?�n&M_wb�hg�"[ٌ�_���P{nt��'�w'��u���	z�|ǲ�np2ؿ]�u�?v���_�� ώ>b>`��Mh����Bϊ��x�j�Y���vh�/%>���AS'�g���	�Q�O�i+ ������������i��_ҿ�1�)��ўO��M!2�{�0��/6��2���{�l�*D�X]+�[��t� �̳�$~6���/�̓�}]A_,]geG��KɌDR8������$��5����Xh�n��5o�2�wR;�����]$+�qHՊ�p��R�B�?c������,H��j��+h�\�����f�����ވ��r�^$�.*�:R�oEk�7��/��8%L��,��"��va��'�W���	� �?q����=�-��x�AG�kLT�,����xD������m@��h-/�W�o�$��Čd�;�V��C�:LC�ZG2���ĳN�0���o ��@��I��	�lx�P�%�e��5�eb��xsN,��y�`�H��mnc��}]�$��)>N.��;��7햧��=�<}J�w�@gh7����� š�^;چ�?�����2��1��
��|I βJ���f�B�QϽ�a��� q�������s�E\�gݰ�t&������z�Y���R���!n5@��FVw�
��y��ءc'C�$r���
��G�#e�/�̤۟���Bè��^�
�a����Vd��Ct�[ßVG2O���P#D�-�sTӴU�rst�^r��h$�<�]����N�#�,
���@�%�%������� �7�G�?[�<(�t��B�����`>%����Z�~|�|�!^��Mp�w׈Z)�������"�����~/9��840�w�}�c����(����X�H\��'Eo�oIТڿ��+��F�d��ȱd�;{�W�_������q�����
�=�
���q�֭Y���3�~B�F�C��lU�q�:����8E�&9�>���:��pB" D�2�TU
m"E��8t5 Kk0�t�`$�ֲR�i�IZ�4*(B�R���݅K�-.QrS��1���z�P!��5� '2��p&B��g�d�Ga2" ����6�F�hw�3v�+T<�g�mk�*/ra(��֠��j���%'u��#|�/�IDX�TB�Z���?��<>�]��vP+�Ϗ&ˈ,��H�so���o�fG׌h/Z4���#_N
�ᦀ��fv�g�_g�9�Fa�L C1@�V�5;��&��^�\�����x�e�=��Cn���,�q��{�5��p5������z��{�ú";�����^�~���#gj��Ji�^㱆��+)���s��3�O�Q�,n��(t��1�pX�|�|)��G׆��Q��O۴��Rl��<� �J5Ar>�ڬ�9_���K7��D��|�O���}�͉�5�i=�iP��=��e�lm�u�L��jw���o�M�d�){g��Q�|�� �$��1��v<�2���f�O�Z+�[g$�bI��VG�{e�ՄBڢe���4�WoMukK�}�tC9]>~�?��|����"(���R73�}(��1'%WApnFC�,���4@si�\�X0"^R�Ġ��]�vd�\��2t�*]�:1'������깏kv�siD����	|¨����'�T�.��
�*UNl"D���"r"�����Sg�"��v�`�<�!V����D�4$b>d����4UƼd+(B���=��;��mx����ݧ�A�nԽ�+��.:�E����Sj�>���ϔ�*��`�+�����lvj-���$N�l���X6������� f�ܥX�Ш���i��D�Y,i2��C�Ɣ�х��[`�Ӈ+Oq��v
pC��.?���?��G� D�Q���:�J�)o�|���\�������9t����\�5���l��]t�j3de�}�.{��U���N↠���|~uF*���)�}M��K�bM�ۈ����!G����h6��~.X����V.
��%h���/��aK������"����2���,�8q����I%�W��x���὞�x����/�XY�0�M)�C�7��io� g\��`J�־s+��<����!��UV5�	'b#=�k\�$�F�ύ���H�oԊl��e��dU~d�[Ә�Erۯ�P{z� ��KǗKm�lj��g�RN�/=�:�0����i6��.
i|9��1~�_:=@��@r>��'7
�^��wkn^}�K���4�;���;������Yg�����[�y{"�;�zų�K���� ?W���MYGz��H�^�N�!��)n��Y!j�R=*;�{���<G���D��j>�JW27!rG����T/��xQ(�U^u��9F���1$:���W:�q���n!�7C#R,Ǔ�M/0@(\%S� �ש^x4�M�&��}��_�d�W�R�&���v����^��qtwt=<eA��.cJa�3�f��l�`& �|���OƏ�?��+��!�ēy`������&����3ރ\[�H���
�@����=t�a�nzY��<de/􇉎G{5f��#�m��i'���)��o���l��C�ςe@�U�#bu!|�̉v�	y���}����&O�t;T˚�<���0p��O���)۽�����'�Ϫ��_�D��j�h�h���I�4��D*�C��ԽHM�e�J'B�>��&d+��W�����J=Ə�/�I>tW�7��T	��i�Y�N��$Ǥ	uٮ�~��fq��|��/X.�e��cR���&�๹�*l�#��m��(�;I����1%[g���llBm�-&n�%���i*�	��hx'W�k���"4e,S�rOQ�M�Ҡ�*ӗZ�U��Ku>2���.��p��'6�H�G��-v&�1���Xk -�C�Jb���Ƅ���`�k�����WM�aj�*P�9�)�(�	9	*k)� q��=>�vZ�T�ά���fF�R��Ԙ��?@���+�.Ϸ�Ԉ��;����xo�Y)���=Fy��̣��Q�1�@R�ߖ�(jsP��eTr�և��-��9�_ꋃ�9?
�)��u��FcDֶ  d\p{��̀(�����d�㗟�ہN�ɀn�vn�!B����ͳQ�����#޾�f� ���'TԢ�1�$%��[�|�������1:d��1�M�<�h4�����t�L��?N�*�ٗ*}�md�����ԋǏ�����q���/��X�&��N����o��� �����_0JVAH��+6���D�������d�ˋ�Z�B�)d��$�q$�h(�c�0����3n���O&k�$p��hyd�u��]�hj8	�N3
3�����b�,�����t�T3���I��*X:�`�jJ6�|,����jJ�����P
ǁK^*t��Ad�\�k$lt9�N�1|7Q�s�L����&��*���p2�j?|i�:��]�U�����9��sG��;z5��� ���pA ar�C�9�I�f4,��h����;��ZO3�;�u���*�&Q��BӗN�� ��&4�-4��D8�v0�T̟��q��H4h{�'rܽa�y��O�'�<\���%���k��e���9�U7x�RT��3iC��&�fgh�Ì��;�Sb�D6!MT)�I�5��Oy�JU*!^ �~����hV�.n5P��\4>A�v��ta�|O��]y��y�q";J
��U����z6���4\�,Im]��oq��NW�1m>��Կ(�]���|�֞�Q���^,˯Tl��'��Uݮ$4���}�E�f���I�f* 2x���O^�����M��婳��vv� ����|���z3���鐅ܷ�.���s*�Z�!7c�"*��yC��D�}(L�Z��Y�J��^>���/h�a)�X��E$�on�����-#��2� 4�Oɣ�� X�����q�d�K�]Bq39@R۷��]/ھ�;���Fí����q�;�#�.`�>q>�8���*��۽�폒�N*��Zn�,�S'&m��ԭ��:���y��������H�U�JeH�?W2z���L9S@\�w��Sf(p��Wqj.ĉ��ET���(�i�a.�H �M�4���&�������Hj�+[Q|��#7S��>7ڀ-%7�^��N�k&!��Rj��+��F�}8zC�q{/�,�������J�|LÚ/5)۟E���bJ~���2�BO�A��y�D�����-�E�*쿂%���j�W�~�g��#�p�Fa�!�'�ּ4{a�kV����L[�B=;�%ݰ-���^� �]h�����&���}mر���NI�[Ms�o��U��e@�j�V�k�;:O��k��:sI�/���Z�,�=n؈�f:4�x�P�+��oNt�U�J�����x��D@�7i��m*�I����"Ds���/.��G
��Lf5Z��|Ih�W
!�1�vk�n ����j̖:rx�.{m���c��]��II9Sr��IX?�iCiѦ�!�2/����>0^p�����7y�4��F?�7L`�p=�y��9�lc���d��k*�G_��j���J��.��xu$N�Э��WFA�P,Bձ� %��ߴ��Tِ��pk�j��K����tv-}#�J�xP(5��Hu�����ex��}������1�,7J���W�7�qaIk�y�����q	
��믨k`O")��[���K*#{��gLH���~Є
C9d���ϊ��]{%�.Yي��.ȫG!N\;�+>27��f��ހM�9VH�	)>�Q\)JN��2..�����{��e|���o�pO��<C�@���I#���/"�/sJƼE�2�����j��z���'jC�$���e���ѥ��[⡲�{&貏q�+#m�K��%�����hJ[�:���s�yy^�cw?DU!��!]ƯI�Z$����P�˜ȓx����UЇ�8���W=�V�q����"NR3_!Ki��leޤ�F�!k�Mt�C�K��[�N�t���a�n]pF�(�_)#V��O�6�Uq�@OF>�n[�!ax��T���X�Dw���bCf4�/�G~=�b�?kNC��+)�T�4�B��{�(��'r��iْp��zrZ����n�"��ݴ�y.�講|�H��]�F�(߾�e�a� #�RMmț!q�����?r�K��:L��W�������϶[��$�/�
��!E!�a.��h-�9:�N,�ʘ�b�����@�q{�Z��c�;��5�5ڡ��W�
���rH�+ld�
�ǙϘ�P+?،;*r��ƥ�ܗ��=�T�&b���]}��ٓy�f�[����6�R�z,���\s��<\�T}{��Q�,�tOS�+?�D6Oy��5�t�
�sz���O�|����l�)��䫒�'�b�Jr�7�g����"}I}i.o`�尋D��IxQ|�q��{�j�j]������[��� �i�y�q��<M�#Xs�j�
�0�Aar�� Y�QN�r���ais����:*B��Z}%�+�=�jo}}A]6x���\����֌s	jӚq>��G.��mh����U|����$����Ph"�T�㷒�P�-FN��ZB6��L��6�⣠j��O��\Y�R]%+@#��� ��̚���:��~b�|���bWyZ�L����t8�����z�؜J4����#6\����z�<:���ź�(���9�t#6d�WE�E�x������,輀��'���U J��Qy�+��n�Iҋ�/ɍ��I��E9�(�r�e��I.  G���6���x����@0%Y+b��Lw]����<,BWd�2�k�*�ݎ:ĮP񛿥���Eֻh��G�2W�� C]�� D��f8*�Y�v0�O��q ��/z�%�E*M�����G��b7̅UH�!���k�a�`����Pv����Kmr1��l-V��5ₙ�~/����m�}�VR\�GS�n�	gz�8=���f�*�--Q.�U'�&����ֳ�9��T��#�< #Ӌb�J���NNL�̕'��������� ���v7�8F�_�p��}<�0&�ŐF�4�>E�+����q�H�Ӷ��E�A�l��ӱӦ>�}�j��?���<�\|	(��"I[�ּ_����T�{��%c j^3�=uT�jX)����"䀴T���%��ڝ�FK�\aYj��G�s>k!��-5A�C��%��'�ǹ !$g�s
��*�u���]�a�
<ꛧ�	:���CP�R&�Ӈ���~:�.�ê��ʒ�NW�2Te�0�_�"I���k ���:�L�$*�'�>u>��c��T�{,���ю�!��x~,HBN���`�F {���ײO8�s�b#�.�o�H�W �D{Y <�|Z��ж
�柁~ԝp��1�3�dnO)����=R_��l+�/R�׾<��0�c�>ҋ��3���=SS9�z��G��OK^�0X��0^��Ǟ�+
zE B:�|�2�1��^j��:��%_Ѫ�4_\˃A��ؘd�@�%�V�L�C&�F!�O%�)Z}�Q�W=�`/`�Bzh��^������$���|�~R���'�G���2�`z��܉ �(>�&=��3.?ƑN�ma!x�B�gg��餀��˦�+��n-�!0B"���n�1PLYz�[~:��+V��K��&G����=)���q����)��Jx���`��)��ǪN^݀kY!c}�v}�wk����V��r2f��"\�H����/�"� U�hCHO�
t���.0�����Ղ����g�l!;�
����`FT�~Ed\��o����g����n����^��(Y�6�='�G����1�.�]��ى�<�MZc#����,m3����L>�`Ui�_oQ��s���������<BIy	["�L
ܜ���_|�w_T������rmh���eG�����gz��3�Np-!+�&�I��Sy4����FvU\��(!�V^hYUA����x_D�Q���pH"($̒��)�/S���gc!�L�>�"�dX�ف����87R���h���.#}�S<���=�Y~�#��g��.�V�ͥ%�iJ �w�զ`��ۿܽ�:�g��E��	�b^&��gp6dQ	�a#ta���i�$�������+��<�(z���W���ϕ#���{�'�p�I�]zIyE�V@��~R}D�@� (���CHؙ��x��������)�|�����Za��U@w���TJ���k�$R.C�0ز���ܬ�rH���T�n�(�,*�+t�6	O�Av��U3�ʰ��=D�
䐃 ��2�	J�@F�� T��Z1��4���|�*S�S3t	s��{�j�0��\�P�y<��]4Z�8Z��
�-<Of��XH�Br��� N�y�1]6z�V�{K�=Ίz�2�O;�U��s��B�����ۦ�®y�:6��Do؟c���
k4�������>��w����<�$��w�*�	;Bz���q��L�y�_�dE1Gd��P����?�����$]��샖q�ӯq;)&\-���m�	9���E%����g/��/|��c:hF�Ftf]��;� [W�?)L�'<9�W��j�������@��$�,O"-��<z���4D֪r߬z���z�JA��U��r2�����SO�5�O4Z�-b��%m� �b�#TI�E�E�tPK��0cp(`P����hu��m��f��j��E�u��Ur����'+,�l���b�t�����~%��R3�����d��,Px
D5km��C��##��6#[
$E-9���%b�1�Uʅ��a��Y�cv���޻-��&��f�H�VK�P��(�O�!��w$qh�𘓫7 �eګ@�d�em ���!3��%}�T�+��|�y����O��x��|�j�:��o֙�̏��Y��&S�а�e�:A9���2Y�2U��?����^u��/�:�Y6�ĭx�g?�|@���Ti���>�I����c[(ʹ�װX��h�io.��GxO�P{�~b�⭕%?N/M�l�6��\��L�p�
{�?���D�w&�%��v>p�?���7$1�$�RIr�����-�W���l���J��A����-����S��*P배�:e�E��r���'	�O�ӇZ�BC�֏U�wc�a�	v=
����Fֲ���ڣn+�ʆk@��$�J���1��&�b 4i g,/�3簣|���A`�o��y8�ex0u  ��b�D����a�45ʃj�\Ah<Θ�������l��8z\l���s��?���(}�2��
��.�h���<���E�G��,=p���w����tџ����I[�;��{s*bZ����� نPҀ��)�'uY�{&>����4�I�ݪ,?�����g�K$�J3B���ѩ�J��Gv��ŢH:���f�7�i��+[�����*J"(0�:�~��#�
������d��>����Κ�DzF��g�N`Ch��<�3֠hY۴q�����<A����:(!!�&�m�l�bKku�Iʽ�>�
�>�mt+�f_u�O�=���[JHK�l���R֥�j�p��pq�'��Ϙ?i�L��9�zls�:��I��z�!�)�Gzct������X��4㸾T�$��_8�E׷�o�Ph󛰳\F:f|.j8���lr@ ����Mf�oI���jJ��`��p�yJ���X��ֶ��t��֚�l�,�� 
܇��e�!k2�[�m�ʀ{c��<�yM���JU|�#���׾>�+Қ�x�s/���,1&��?
Q%��QD&��m�^(뵕����=�B��C�|��ܒ�mM��z �$�hIE3Z'��I���s���L���ЋB�����`�!�]�_���Ȓ���ʧ��y����>G�tr�� �؇�F��
�2�0����{�~¸G[�.2�CGa�\��1�,ig�FOY8ޱ����y�K����(0��D�`�]ïV�egZ�>��Eجh0�cf9K"�^������&H��	9+�"��?���J }"y�uf�F�gPg7��N���T`��R[�Tk�!�"�ҵh�Wa��s\�s*u}�m���X�7�1�dw��4�r@5 �� ��@��#�sK��7R曝�.oK������;G��H�fe(٫���l?44��I�SD��)�Ǽ������3������c�K�Բa6�N$e�)�r/Zl!p��aw�
.��~3�VK�t+.A ���x�gU����:�~��l�tb�=@@8c,�z�E��-W'�eg���n�{��UCL59@W%4������ᖔ�Y�����O`"�l(]U<B��(��/���͞�-ǵ�[�Ĝq����3Y�� �k_F��0�&�^h:�̒o����˫��ᑦ����l �+�3!���0�5�`hv�z�	4S&��o�~�N������n��
%¦��ʒWb�r�Ramsv��mϦ��3�*�$��y��~�EpH����`@�����h��*Lj�����R^�6�E�+>��+��DtjG�;_ό
��"ZU:ݝ��[Ps������ux҈f�
�x!�Z����Q#���(�I7�G�o�{CQCA�T՝r�����P��m��7E���|����ڤdV�6u�̡\#4��Ն�,'��*��U���ߧ\�a��u��'zDKQd.l�;����K��pY���K.�MH��غ$�ח&�s��w�J�I�Z�u�QI�\:]u���v�3!u"�G��6��
!�^��Y�#�v�}�I0���A�+���R��ne�2�J���Jy^ts�|J�[FA�c�a��c' ��n~�b�e4Ck<Ys-V����ZeF>�;�<�nH/�4�)�hH��)߈��*.�0;����l�Z@u�z�b��í�4��w0�k��$��I��/�Z����pl�-�Ԗ^�|��KU�|���^A��^ïs���:Y`�_�<ز�&^����^D���r��;�%��ಹ�a:H����G��u��iHQ��8+���(0��2��At(�����oIE�b@Ϩ/�!���>�0�M�){����c��q���NH�m�x�!�P/n�N?R&�z�|�hd�3�^5$[L�[zQEU �nM� ��D�*���	;4ju�t�9kV�[ ^qmc���_��B������7��}6��r��숽h�'�>��U�h�]���y�%�BH��T��8QuTϢn�N��liF����\��y�aگ����^�&�80����ֳ�T�?%m�>��5�������2�^�7=ς4��ޫ�)���U�H�e.dz��~=̗:��+����g>8��̤4L� �_�k��Z�,�|�X�A��zw*�a��m�xo�R���d���&h����m� $��?Gd xɚ���.zK���<j`�)�+�ݬ�Q��ڊUaό�:|\��V=%FCW���v~���'��1�����c*Q��ǲ��l~^��TI`6�o���L��q�9s�ʷ��}^�n������5���2�?�|�OL�D�uC
� /Μ�0Ǉ�T@���ƹ���I|�)TY_-�����[%o�9��NB#��6��Y	�J5Z ���d����3�r�lU	��9D� ��㧝��|������+�{s��U�*c~�e�Q)!+d�6���z�N#�Kx ؗw%5�ʀ�Z#�+�f�/�he��9�v�o�V[0CGg��q����K�4�}#)�Ǧ�l�1�.f��� ��F&/�m���yeU�U��C�,�w�c����H_K2�& �s���D&�`��ץ�5 �|�>��xKX�"G����p�Ծ�tOkG�b_^�	ӽ=n��%*`-xA�S��5ߊ�� J��y-~���
-E�UT{�Ӭ(N4���E���r�T����y|�����(�5���kt�U�vv�McGIT1��ݴ]S��Ú�iS#��/_�K�)-��hb".�t���VB]`�&��DL� �f����2�:��<n�[�aR2q�C��h�JS}Gҳ%1J�2�J0�¬>bJ�����n>�ԔΗ���p.�c�����c;Ҥ� �{*Y[Ϸ�bU��^�(��}��5M��q�"��S2n�(��!�E�3��u5�X����
j�Zf��S5�L�9`nS5!	AH����yM�wjfcځ�V ����n>C����m�2��Q5��ݵ��+�Z���zcЩ#D�_n4p�pvQ������E�f��A�\I�'���V�#:����D���\a@���0�pOR�)ڝ��G���3��]�ϔ�cq/*�9y��(�����e�2��&��79���ul.���%6�x�.Wɹ�Y|.�����թ+{�1b�.!�]qV5�Q�7 p�0��͎̓	���w4�cm��Į�!ע�|1�g���|�H�1�n�����N�E����{���/K^O2G������}&oL�F���C~^�xߓҏ�2͂�2�(uH=85�gT���W�����چ�ۖ����Uz�~������!�t���7����9�?a�ޯH��+�����HIÈ����or�����*�x��Y6ќ�$Zz~_�E7Fj*ߦ�&잨��Ƀ9��8�  {��9�{*���iL4_�X���� �����=���<��0�HE)��Z��h�@ܾ)Ť�e��.�<@�u�(�&�&tzx�a��C�[zص��1wh���� S��j�|���|	�	V*�����=_��yԂ���yɔ����#�n��S��4�;�;��U��o�oQx1тK��	��~�W��y����O��$NQZ-(�u���`ߟށ�����>IFU�u g%+��acX�K�b�f� N��I F.t��[�� �gy�v߆6�h��朠�`#�؍��f|�LALJ&T���k��a��
*��z�YM"�G��@7�|T�x�s�
�����<�m����p��?Լ���C�����L?�7����6��i]�XZ)���riڡޙ�A�`+X�bcǲǜi¢\�y8�n����2د�/~Xc���ݸ�.t�~�F�9;�&V�n�����������/h�A�L�>�$1�j��d���J����48�6v�0�Rt��n'����5M�#��`᩻	b8x��,��65�����dHeeV�:1��X^7�_.خ��eJe3=bx��yq�ʌu ���W���cP�괟SӅ����A(-Vr���Í����>[�I\�����}	�2��c��O��@:�m�V���'}��ɉ\���&4EI�Zk��*V�5>�D/���ŭ�Շ(�
��kt7^��L�rj�S�ɱ�YfjS�zc��%�0(���|	�8���$�t�}<���Z�-O�p�`o{V���ƒG����8���qT��4�Zj�ƨ�50)�^T6�4�8��9�R�3��y �T�����0�L�p�m�p�z���a���e�K���"G@��+r3zi�I��Q�ly7��a��� �
�&�t&��,�)J��7��GU*{�ӌ_�l��b�홖O�1ߧ���R�O0���<�����X��5�������x�\�fB�kb~�*�Vy�>�~�?�1g�$�c�f<���.@w��"@G���`G���P�^ۧ�آ3&��Ft9]-��
P���U��v��*�k7����_}�	4�|qX�O��˵`�:�<��À�7Ɋ��B��E��f*`$@C�gB����KjX���WU��
�j��Y�g��쒲�6靖GgGų�k�̤'���һ��tȍIB�8�VF^
Q���u����Y�7�V�CB�K�&ϖ�#,��f�����,���g����n7	��C�i�义!`b�S,�n�ul�/��ƌ�H��0���L <5���}r�`�u�v��h��un���`WP�5c��58N��R�#�&��A���j�ʣ�u
s�+���߿�[2�7%SJ����nю��qŨi[m���J�h�r�t�����pZ��Y���ȞXF����6.���KE>�$�7vK_���#I��Uf��s�t8��M+)^΋ņhc�sy��S�!g���3���S&CL�e�F�����I���p�ߙ3Ui.ۥ�}�/T�RI+��������� ��k�����T�
,�8�/�|��k}-;�Jݝ��L��������k
j�ըb�����*�5C�q���p�!n�~s�驲��ke]���C�xhm�V��d��z�5�|�O
?��䐞�|���]�"�
:7����!��rJ��j�(5b��ٖg� ,���_�<ɖkI'Q%�3�1VA9R�X�^�X�W�3��N� ��dÕ���jI�� �X~*4y8������섌};w�y�[����Ϲd�^H5R��w]�~�r6���^��T[ ��P�֨�/JO���V�oB�cG'�_��:,�j���y8g+�_
�g9��.�������X��bj����;"�cJw�h��5�߻��'�����6��cl_䭌���]E�
gn�$����։�d�f���c#�k-�I���L	L!��W�4e��h{�����w�����.~���Xux����=D�Riшƽ�]{D�1�^�E�Ǎ>[���m��k!K��#�8�wȿfZKr0�La}���z�Ȩ��c���4�L��3m��p���e]�;��:�F�耓�{3xDĿk[<i�~|3<1� �\G�i�*`%�"^��2(��2a�s��OT���g���,���.h7��9Qgf9Y�
7��M�I�Fa��E��7����f��Yz�8�� ��� {i���y�!P��&a3
L�CK:8n���������~$a(���:�}A�5cm<ش��"#�U�$��2�F�V�EQ��w@d��耦�(�^��P�WX�!���
۬�%�^v��dÔ�s\���Q�>�|����U��~�-�3E`O32�@ng ����,8�O�Bmc���FB�g���=�(Y�̉�Qtx��_q�6 L;�S:ݽ��g���h�Eb�.�n�{����]�H3��|�+��5���z�3 j������!(��O��䰴-kW�//@��@�E;����$z�ү
��*]�H@2z�+P������3��g�������%���Q���� �r�1)k]6;@�Ւ�vbl�[�Vu7���R��r��!e�A���B%Y���Ry�oF0�9>�����(>=y�	�_�[��-aL�Cn�)�� s�t��Nt�2����#��N������/]S�.�|�{�k�|�Ӗ�w�+�xЊ#%�@5�:���O�Q~4@ߣ�� Z�Y�r���T��1{%� �z�)"k/����u�آv�cKl�E5���=�^J�H3a�¶(�����zNSU��,v������մ:�G]��w�F�{g�]�˫r�2���%҄$u�=qHwH?h��q���n5\��:'d��g�e�'(n�T�h6vai!������a���b	�Ɯ9���o`j�x'�L�8?�� �I�3�.^S����p��4�k�S�%�Y�@N�!y0D�y���F�!a��3,&侾���v-C�*u�'o��� Q1�kK�t�8�m��elbw\�" �sA`�%Y��R���ޥ��;@;�8#�΅/^OiH�Q,^����4H�>�Z�U2x�A�k8�
Z"��ko:�H��BF� Qp+w�V��/MUT�A;�~�S�^FM�8�x��y����
0 ��:��:����>��N����c#Fb,7%P�-�ǵ�������l�p�_����`t���]U	P��HY'%(�W����Vo�r(�;c9w¹3|���>v���8�1�}դksk8��-�I�����ɢ���3د��㖏\xq?�N'��f�$D?1�hdw��C���t�8~
+&�d�k%Js�����~��w���b�)2������'�|Y"e�^D6����:ls|/fO�TQ9c�����%����w�o�k�B�:؁���N5��7u���UT;s�$��~4:^d�����M�4��U6q�L@����V�X5׎�UƊ�]��6A��2S�e�*��=8�����9��McQ���kA�����?�C_����h;�*����ƫ�Fj������j֟I���y$,7[{���s��^���� ��{�O�z
�~Z��:h�����	g?�T���n���w��j��h��@���>`a���&M��<�3���/�Օr^�4:b��EǨS� �V���8�'M�d��XP�8YťE,7����^aw8�C���a�L��a�P�㙽�v\\ ��L�L�D����'�q\J&$*Fa� ֐���Ґ_|H.�(Q�tɬ����+�1ɭ�#���JUd	��~"]�u���.	3K��J#���5�f�LP�f>�>'V��;3}� <�@�_�=|R^2E��[��«��0
�"L}Z0����a��|^V�	1@������̆e���W&
wQ���>�ŀ֣~	P��!�?[�V�*# ����A�1S}���թ��hrm��7�f�L���Hr��=�w� �9��*�X���H^ߗ��4��[b��k�#Ge-�'|�/B��}:�$m�{��)���i���i�t�,��&Û����h��v;����m.K�n9iz�
dB�E��ʐ�HA4Q]����ӛ1��>Ɖo�K$dm����l��B{�o��W��$���n~���g����ˁ7��->9��4�U��ˌ�;��Q����cݪ:�R�t�G�r��I.Y�j��?ğ��~;t�$H:�'��[�`M�D��1]L&.o�3t��Iå�Eٕ��}�ke���-���yNǃȯV�g���=�Pڄ��U5E�������99��"���t��L�b�g����G&X|��yFA��ƇY�d���o�N,E�e�� �u"��������,;i�b���N�	�z�m��"6�<>GL��sI��0�s��&b`l���D��H�߾S�����f2p�`���l� B���}w
K�87)h'!�N�8U�J#��e�Zw� _ ���
��J�[3�c�o*�믑�P�fdv�����s�e#y|o�_�~HO���u��E��Kz��<�:�����#1��ߡBT�谰�фWOOq�F��52�FpjG&�)P9�Y��	(�lE��6��c{4PK� hӣ��U��x5QS�X��]�n�+[�fb��L�ދ�[��%�:t���۬^���`/��xonռ�ܬZ4	o�.���5�c�R��e�q�G[_�Up�g-�����U�qFM�$9er L�Y̾�Ee�Z�����P��N�}e�+0��>y<z["ɀƢ��J�@��ޕ�C�=��⟸Z�Q_�qҲ5T�#|y��>� ��g]��o���:��E�$��B�_[zgͪ�2��H:&�©�Y;J��+_�ڦ:���D$�n쥿(��>�vQ�,�'�G�^y
Z0�����g`�&	��_������.�p�AC����WRE3�� ��Kwng���?rEzok��W���dڵ�0+�ˠa�,��O�:A'� �������2�2*`hS� i hte��)���"��6�ޏ�h�兖#���6��G��lL/1u'�V�Z��������?�2;�'q-a����@z���s �|���쮓�����#��c��T��N��CbF�&�_(
����ͦ�u��9��l�-}�H@|[(Eέ�X���I"���"�eJGS;�yDlc�&�YOSx-ƮӜ�I����o�$h��nHdr\^��}ܸ��͖V��W�	UU{���E������������r�w��`��cճ�[�����U��M�"p2�2��V*�fY?A'��:��T�e���� X f�3B6Z��aV��﷖��f��,� ��:TΉ��I���� s�a�Mb΅��[��d&v�_�f���KE�4 ����fؼ�w*
�U��v]�14� >�W�W��'�6�ll��n���L�M�����$�%�b�������2���\=?�ۙ��)��
��Rf���Ub��ߩ��`[W������02ZW}r�K��eⴕt#Ԇbl.OԺt,&�#��Y6�6©��7��j�i�,���k�������ct��!�q���ew8�(��Ef�H]z	���h�@c���ա#<�]��+����ͱ#�Y��xK£�W
ԈM�V�Eup��٤��cM����Щ�)Ny�]�29lF/Je��l,������_�B@3$��Ļ��,XG�N#�ەX�;��Dx�~�����w��7#��u��}#��Y�A���Q?��$����&� �)#ar?�`��U�1H�]�J�$vp`��EQ��̴��i��,�ӟ�OQ���t�X{�b�sG�Y�w�B3}t��y-Ҩ�"���rƥ��uD�&��#Wy�u>�
߬5��=��\��T�E`����iD"J� <��X|J))�3�O;��:��ܻ�+�y���,V�:���%�V����s&޲�;&�v��\:�?R����-�K�V�Y}aE��X�8��3D�WiKI�1���K{�"c����V���v�nЀ��_dr�?lm���@)f��)_�P'4	�bg~�S�b�J�oM��n�ƪ��ڳ�q���Y�/���B3�yS"����>�I3Nj"K���YƤ������zJk�u�jPy㴊U�LU�{��6�?JP9@�ž�K�~Ǘ����ݑO����Ou��i}~��pOF%j���Ǝ���j����
IIN�W�uqK���O�՝qy�3؊�h��^��5)0�V:�Y�=3�3,��&H1?%9��dnƷ~E!�����qO1I�{	�w��Q(����<H�y`Š&'��J܄�"��_�ӆ����^��6. ���J���=!|[��4�kO�ۛ_��-&�x� f�#:j��F:�0�}<O�a�e>�����#��Z�*��Nă�< �2��f~$>_��o��H���O髟��<�/b�I���TH����Z��H�B�?>�=�=�����O78��{�}uns�Z�}�NL��g�\/:�/��)ŀ��H�7�y�HI�+w+�mf�D��f��t곽�`�i�vMGg���f�YC�6c���l��?C��jmo���� 8�L��e�*nl���_����6�Ex~���+�����Z<�����>(to1��?�^�p�V�Ї��F�Wl�����x����%�4d���h��:���F�^�[��1CuX����B-��������/&�Rza���r�����(���������|l�h�=vNE^X�����E3����iH\4���g�n�}'�(v}!�ࠌ֍0��U���sT~]L�`�4�W)�s$��`B�!\�t6��]&M�����,]:u6�7 ����3��i�qd��Od��+Zc�ė�,~
��HUs���{��b�۬VI{9�;�j�t�Ŋ�|A��F6P+W�T���
�f$1	����'n�O/ź��pV�&*\�[�����B1�O�K@u䓠Y��Մ�m�q�:�c �_�`⾮)����KMҠ���E�V�It$����؈|�����10�?Ҁ;�I�)Vl��Fkr�����Ѕ�W�L�6��˽�r�<U�Qr����X,eQ�8���POe�YnͶu ��F��\�\w+:9ا��%n�m��.>w�Xm��1�탂+ ��ʣ�8hu��,@� t�H���P}Fu��ˈ=�	�H�����Wg�f���sb�F��n� �N`�B�= eG���D�􈊅��+��i�>�|�O�&�Ȕ����zd):#zD�et�9�&Xm���x�� ��q�>q�.nǯu�#�hq��7x�${5<��$���_�o!�ֿ!3gF�Q�m�����H 4ل]d��	4�w!FZx����b����fu�WI�o:��l���=�A�7�яC��+p1"R��Ά=GP!�v���q �������:+iPa�]�Ǿ�?��7u.�=VH������Ta��3�!ƾ�Vd2���qT�%�B��;��i��b��\�9F�W�ѵ��s�0p�h�b�/,:ڣ�<�������[���5�(�Zׅ��0���!�\�j*�5����"0Tk�A�5�]U��4٠��20+O����tFۼ\�*|��ц[,�f�v%_��H�#S��s%�������YqR)�*+DѓT�VU@�H6�)���C�̀4�$�
�����2|�^��[u{�����D��@�D�?{�15�֣n1��Z��=���(���f>���0�Q��l�5�E�3�����ewd�n��W�+��s�C<u�pW�&���8���P�̻����;T�KlsrI$�r�?)�����5bR�Urh�T �B'd�%��,ӭD</���0^:�ӝ�q�FT�;�^��F��D�sC�/��@�#]�u ~�s �{"���1��P�K�B�l$lFG�FR�u��עF`8>v9�T�)��_��Iq.�Be�1?��=�m�/oL�
S��@�4|�T,}���ҡt�O�?&p���[$�d�[��n�%2	�ET�U�&ηk,g�%*��q:�����D�| 4|h�<�BT������zt��{D﵋FUj��� q�����a�G^�8n@ ���Wq�W��:���{�Mf���2u"c14�)��']l�)l�m��$S�|�;Ј���\�x��
�L2*R���MF8n�3�˂	!5�6=����s[
.c��� �ѻѤ�9?,-d��l]��^�B4tѳ�˪�\�s`������OB<}*v�D�H���GN4�.@������E���#�D~��Z���E!�t_ �NY�:�˜���/)�B*�bԸ�����zU���p�x�s/���mK~�<O�D�����ڎX��Ļ+�H;fv�����@�V����	k�<;��e�RE�
��X"��];Ӹ�9"���7Qy��}�2A.>��V&e}�.���6��ň}&p��L�� `� �X�#^85��u̫�Y"�2��@�@ ,h2c�Ω�W�Zɹ��A,��	?wK��)�^����ֵ#&�&�[�/�����|�A^�r_�#��j��������k3_0~��C��2̈́n0C�𴓵V숡���oC���iffzSݡ<Z>������XIѻ`xߝ�j'�E,0Gp�;�]��顏 �]��Q�E�yP޷*�XF�Ky�g
Ltuw!P�ۃMiI�6*�j"�������v��.+�K�А��[�x�f(J��������U���56g�a��Ѵ��JK�0$A�]f?��*2�B 1�zJ��a�{mL���t���Hx��Ep��;P��vǻ��Ia�QhDp$;�G�o�Y��3y[O���c|ƨE6�
� �.�㊎���H?�H�Uot���0--*Z����m�7}|�w�h^_��|�����< v�*���&�8q�`�w�bʠ.�(�~��_9��򎌸�#�Q���rә�����I���&����W��(.�XK�=s��^�qfZ��.il�9�ol�Ugv�NU����Ǚټ�6=�F��6ns���;j��g�ψk���m�m9>��N����C��n���{=�Z%�t�S��?��}���_�B]6�j-��?aM�C�^������\}���,sM����5�6�3 @v����_<X?@��d�; /!���W,�/Fo�e�t{�m���'}RI�KoD���_wD�n�[�ջ�	��%����+��
p]��q���C���>������d3�ҁ=�/L�[��6��,���5�K��귒i�>j!�M�c_1�|z��C�Ҁ������RT�'/2V��>�ȰU��{B��[��L��_B���ZCѺ�N�l�~�����*#Ĩ����b��`���m�V��蕽6�l�Jo��A]�2�RZІu��s͡�/�u�C��ǩ�	Y�A�����	���m`��=aj}i�'��� Ѓ�N:�cz�4< �v�}���J����^���?Ս��<^�������nX���@UT���լ�(c'y��B��.#�$7��"��|��F�Y]>°LM|9I]�D�C��d=����2�?��Z�tjs)�������������ύѥY�$� !lcUf��%R�������|��s���]�J�{��ÓJ�la���P_��p*�0!ہ�i��X��P��EFA�v&t����kĭWZ\���O��Q��}Vaz[��B>��$�"�a�e����[,�j޹w|*N8�gǑ�`��`��4�1�+�_��|����j��["tޯ��_D-#��)�S�8of�����Q�x���v�<�mQ��֩��@k���RE�^k4�9ɤ���<["���9�)��C�~G��.�-�خ5#���z���]�y�#S+�����d雅�i]=��q��piV�o�z[e<�<�p����
�F�\��݈r�H�)�Z���߈�*�%So�[LF��i��Z�_�=r�'�"k�gF~K%�c�K~�C\���R�l����;�(0@z��ez3�&���c�a�`�b�E �ꏨ7���ߙ��������VA��i��?��\R�R��yD!\��c�ϼY�pk}#G���hjɠU���ނ�ax���;����(o}��G"	����ş���Im���?C ��똻v;�^۶連MJ���u��|Bye��/�P�F����z̈́O |�i�0�����ʺn��ߴ�)t��"*�/J���ǥ�%X{Q3;)�W�R��B�O$��&{��]�
�t_�M���k�+�xUۡyd�t;ZR�Iq%��J�^�U����Y���=�$u)FGuZOT��rUěT	~s��gr_�%��"�q>�e�e�oƜY��zK�ϭd`�i�_��SٶD~�NIT ӡf>��˳|�+��.놋w�"$����;��v _���_���BkN�^lFEֻ���I�/ܞ����f�l�-���$C�������Zf�̂���؎97g��׉�g>�K%���jA���Hy>�X��(5���oK����h�g��$�����8�v ������=����}�h��$�.8�� g�/�Ϛ�E����L�J���p�Pw���V��g�0�?��
��X�F��?Uq���p�w�΢�O��IC$${~ٟ�3������-k<ξI��VN<���a�[�%-
l}y�E����������ѿ'��y��u&�j��av���5���ra�;�ύY/�!a��7�O��Gt������+&�ƶE{V���Lv�IsY�Ҭ~��;~��pNb�L�9���&m�T��C��q�'�ĳ,�hq1�y�����\Ĉޏ�s*+&��T��^��s��1�'�j#�XN�\R��~��R��3��.�bp��U�P����4��F3]��Pȍ-���go�(���S�b������>�cj5�%�� ��-��A%`S�0*޼��^�$����_�dJ�";�m�EdJ�\gH0r�Ĩz�/G .F�����%�j�ZBf�`���~%���?�B_�"Fn��g�s%�9Z��*6�VKy��*�����Td�}�a>n��^��Y�6�ۤ��?��a�P	�AF�\��W7�\~�}|���u��Y�\mc�����[��ge���o�������d��0�����r���Z]�}�G[&z����QO^c`�@3K����{��ܐ;6[�$�&�{G���+)w�U�g��K&������iU�gx?���sVQ`�0񽃚J�r�
xP�f�-d��k_V�8;X{�f�НcNL���U����$�O�������k�ܱ��9j7�mc���tT��B��f$�C�'�	����ʌ��M8�L\����R�p8e]P��}�Őbr��h�ŕ*3UȺ�X��=��,[m�"0@#��!��a��^<&L��D7���<�+ݵ[f�����ע-ؠ�L��c���V6���=�,������-�Yq�Y�� ��B���&�N)�e�_�3
�����i�`��н�I�HI��a�n�3*�|��z8 4Çj���GO����Z�*t�����~ h:�� "�5��&�2�a��ơ�8WϘ�ޟ-�s�d��-o�V#,�	T�Y2���-С U���9:{�C�D���t�Z�:O���Ziat��z�-�̓{	�*j�����]��(!~E&������3K���M=�4�K�VM��j��Պ���gU +�]��a�{O�p�#M����B�2���'���CLg��Ѐ2�d&4=\�r������y���;Ū�ǃ����yV��������U��-))��$y̘>;�	� in��R惪�F���S�iK<a�W��`���u)X��Jߎ�(�}n��Vrf` n�d�˧L��4j��G�R*/v��q6�Ϩhg��hF�_�e4ҽ.[d�˄A�&��n��;�����:��YW�L_��x��D-�����K=��*<&�?�+.�`���ì���o�ߨ�s)�n�Fm&��BR�z��ڄJ �Y�� Y�|y��9�
Y�#e���A$ε&S�Jn�4�x��[�M�z�E҉�_S�X��%�q���ƪ��/c���uj��H�7��5-J6V{<��ਙ�E&/�H��������u`�l� 5P\��B��4h^�p#Є$�C���G�ؿ؄��v��XR�����Pl���d��S��b�w�����O�.K)���	����Y	[�)��6y��o���S���W�$�%Xh��/	{�ƀ��+�����)+P���ѱ��: ��[�k������~^�:���b�t�`�r�xvbh��A�� ���!�un�6V�jhš'��U�<ؿnf����&}����tU���ޖP�ww�xLW��t͞,[�!�:);��<�m�<�:�O�j�u���#I��uJ�f/Q5�Ƚ�Y�	�������${+�ؾ6k�2S��[���p�D��~Ր�S�c|K�� 6�PA�_�H2�*��8�`:z�ļ�/fϑ'�[1�r�M?�r�$�ZZ�ŠO�96���ݐ�_������ݬ���Q���8Z��H��Ҥ(ݒ����f�筘�[dl��~�c8M��i�fh��*�#s�QmcM������	���e�P��˭�;̺]��E?a쌢��S��+�/��ο�'?T*/��+?pX���R���G������g���5xӼׂ��4�ī���  ���'2T~b�ِR�f�lC�3��dlTh�x3�Y9�q���tk���ZY*���D������2�à4�S���J��`	R#'tM��KkN�ͳ��rX�[���Wq:�|��u�soI���ٍ�K� MM}���䩂�c)dgB[n9dE.��������Ϳ�������$�����@ǜ�Xq��BN��u���-(Uk�fV����NU쫖��>��R����e��Y�:h$U�f��E0�4$]�ޒ�� ��c�	J�+ԑK�?� ͡�bo���*CWCM�B~����>��HW|Z7D+BA�$~�±���,b�m�[�կ
ć��+?�k��\��ɠ�v,\����H��(�/Te�Pf<����R��.��E���Jecl,󆇕�U���TNվ��a�Nm�ӟk,D	� ���T�[�L�>��t���.rӓ�\Q2i����:2��(L��̕̩��s�y��MhGmXx�*��9G4r7ѳ0TtH���v�x'ϼ������?�nħ�6��7,gb�A�	�	�����)Z>��s����9�a��6�U�0��������/���	���q�w<U�0�glz��e�S��|jF�h�Y
���W�E�GZ�u�a��1a���˹ih�*ƈ�R���/
q�uǐ�(�Udu���0ܔ� .��AR�y���K�R!�H�=dt�xj�V��Xz�B䵌eg��MxRi:姍�E=zj��.4���4��䂴���;X�*�N� �U� �F�7���F��^��+��RO��Km��[�6 �\�[5��/Q@S0��)�8%����P$H�C�׮�&xb<]�<E�r�ǔӜPz�w����,v�(���8UuS
#d`"�W>����H2R=�̘�e��.PT�3��W���X\����G�w���0�@%U�p/�?�_i���w�و~��{z.E�����5��	/]ߺ���ڪ���¬ml��m�k�Q:[��6TȾ$V&+Eg� ˓����C����,.J��O�����_���S}�CK�Y�C����2Yu�ؗ@�qd�7���8y6�
�dRߗ�p����ɪk������~�J/H �GOŴ�ҔCd=B�n1K�^7�-�5�}Yw	7ʳ赬c�'?~�JԈ}�}v�����(���d�Km�}hP(y	�}��	�_nS#M��#�v��]���0���"���'��\�M��a|�@�f�N�IB���f��~���p3����H�Roy��MFk�S���ɿ?��2�L��i��`-ˌR����#`��@� ��W|z���B�4&�V,0���-�b�<����[8��V�IΘ;1�������/خ�ng�D��m\[�ǽzRd~s.2Hۿ	����=%q �ێI�}x��Y��#��Y��c�0�ȡǗ��E����M�Q>�C�����n��,��ͪ���Ff���ۊ�t�b�.�F�0�k���3E���_\=�}E�Hg��Ka1�kb�	�MQ������9���Ĭk_ȳ���i�xJ����M�[jb,����}^���ܦ�����GB<*C��*�����6h��Z���aNk)�O�VK����:���8�.��Ad�j�G����.�Y�m5:�`�35�%Z�xM�O��m���wm|�V����n@�|vs|���b���$��\�����֪��³�7J.��S���-��_��QdTw3��V߽�;��A-��<;���wP�O�	A��]
�U |=��1q[��L��=��aK�A��!轳�����N����V�٥��4y)��<j|l���>���SK'\���EN��F�UȌ�qd*���NZ�%�k4\O×Y����;*V8|ߤN"c�sA�˧����3�f��N��cT :r!���w��.��D�Ɠ����̓a50ؘ)��z����w_L�UpZ���B����qj�MI���b�u�/x ��c��"�n�VQ�+��M��!S�|�eze��S;{�O�Zu3��t��"��G#�����j�ҿ������c�HT�}�O#U�j���E;x)��g�����l��+��-Δ �9t����;ϒ���,���r�$��3�.�p�ڂ�����,_yb2�H�6ۼB\�#��	k��Q2qM���׳�'����RG�����xD�1���Ѓ�1>>����50 �s��WsV#����p&4��hWg"N�A�w ��*�+'F^ڔ@j���w���Ȕ��$�[�_��&vj�o8/Tq_�}ub��o������`��q����{f!��G-a���GF����
���S�WF�w�q6xe�[�5����J�E�{�ؐJT.��2�,)9����tp�j C��pĚTD0I�.�#��2���&�����^���n�K�`�����24���JҒ�ʢ�����Q?�6e!���i�at�6��1�(n4%(,`Y�׿
_Sf�'�|�~١�����n�Ҏ��Η �����N�Z�E)XO��- �,��*�~�E��BC�oZ5�,ܧF��Z��5�������>h�$�93�e-z�5�@�r���$@����F4
nAw5qv��W���	�7������bIL�����-dO�-b�Yl��U�F������Mh�3�鈐c��K���6a��~���i���j��i�n��������ԫ�>N1�-���l����ɚͿh�h�����`�oB���ޣF��������uPBP����I4%�s����k%��A�s�����z�Y��~�co��\��y5�B�B���HXѶ��~��<�����=Z�{���S��06�*"f��o[CǊ���Ӯ��)����Ř�X��� ]�T��z����U�B�C�$�d�[��wiiFx�^�E U�M�YJXӦ��[SV�'�/��H�X���8]2EϺ�<�w{L��\��;���䕏>3P�����e���������g�ٰa o�&�<�ʾ�e�jF���`e���ՔrZ2���-���Z�m��G[_w���t��7r���W�4t:f�4o��\0�%I͒["��;Jǒ/�*	4f����,�:I�~�PӢ��ޭ���V=���f�zr}4�"�ﯶ	6���qyg��a�Y�����u���8��S���鎭�v�~@;I��,����}`VC_eUUm��kl8���$m{!;p��	ී	��d8;H����)\y����3z�w����f��i�쇭+�G�[���oQ`��ONZ��������~��.	�XMP���ͯ`[A<�:lG��"TT��`�~�q�H`��wX�^��W�[l���Ѻj����������A�n#I~��0IĄ7��gv<͡�rŊ��eFġ`yd=�H\�bp�]��<w�sp�sddb����rJ��ۋ|�#<f&�w��_'�^�%�P6��i�z�ڦ�>�g���ܻ���2�����RE���(v�(�cs�/F}�=Ǣ�[���	x���c$�~�e�I``L����P+�(����<���:�Y�'��Q7�#�a[����,�	�%K��L��+%�� ,m��f� 	���V�#�î�mX�����Ω�
�x�-�}
����G�����,�xO�\ۻ�גo��"��l�]�2r��b��Τ�lF�O�_)�VV���@�dJ���T�^� o��|���5x'"A��lL\[��|V��@<�+��xC&09RT�����9@3I��Z�;حզ�5���A�'�T�5�4�!��xK�K�.VA�X�b��;y�P�eˈ?�R�13��76}#��+=u��PjZ�)%B�)�L�h=a�~߶Rj�6!
��[6����P?Щ�^_G[��ؽ�-5���i���w5�2V(�
s	Dt�?k.Jb|R�a�?l�����ε�%�&�X�wVKu*�C�k'bc/Dy�}����$��T �I���9���2\� e�F��c�>��������UG<�f��ߣ5*�|��Fix�ψJ��Z>|��=Ĉ�'�3;�p�������c�ƴH~�ԸS<��o
s$�&�`=��"~��ά�k.�8��ʚ%w��`Qr����-΄d�a�u?�j�ᘗ�5���e���-c&���[�6�k��T��$��K1�'=�B�tԠ�JZQ�w<���N^�9x�]�)� 1��;��@�zB�qSK�s�%��u�4�g4�a��L�il���w8�p*W� yy���y��|2�0��x�LbMgd�B���yL[m�̣@��@:,����){���	�S���,p����~)��Hw=1��:���Nt�Y�.f`��쬹���o���:8	�b�&���P���<�����ˮ����k�9�m6�C��ލj�Lz>;����bc�	a*p��p�7t�.+P/A�3�mkr�RYۙ�V��0��U�+(l��)�%�m�&��L{qʪ�)���W�����x��b%� a���!���I�������D����������xb,����"W"��:h�A�I���=|��\Rqڛ�>����*+�j�,?_�~��hJ|��s���WB"���,%���I���yUB|�h�,ؤ0�0d�jkX*3�����	2A���K�9�	���1��6P.ԏ���v�Z1�K�ue�9�&�Zܦ�*)7bg�9���ZXFh"z�`�X��QsBj$��f�2�. B��&cr��W�hS�?Y9�ׄ��;Ք*ӲK,�ŏݫ(|�@�U;� �?v7w�~�(�de=�o5eα�c�q�ʔ$%��?�/�����U� }3�&7�H�ކ����[��^ ��e��2wj%�����Wp<���e �H|d�_V)϶��[@�w����z�3Ē4�# Ee����O���e�.Ù��Ў���g�5� �	���$�)��Ԯs�dv��������p���}���q�Lvk<Q Zk���� ��Z��S���uKh�E�� f���M遞����/�̄ ��+3��c�f���'@�ЖF�1��3�Y�u*�EkE��S�����k�Q-��y�V2���D��x���Pw��l���֌ �x����I0�y�<�%3��;Z��|E��$˘��	�$YO}n
��(���>�Y�d���4Zc�㪡�=����h�)KN�7�c����[^�xT��0��_���\��o4�V'��zW�p�ʳ�篤�%P�O�z��p�����ނ'	�/�2���/�k�_�J��)��Tk���N|3��J0Ͱ~��뤓�ʬ����U
dlI5m`x���~)�N��UΥG!Q�_�x�:s��Ϛ��.v�aͷ�tF��9LY�lmg����?  �p���L�7�<����e5W�̧6��R'z��6�hW��o��#�Dk5�� �{ء�R��ŗI���V؅��Ȓ����5����[@|��R?˚�k�P<jD���_k�v7�� �w�00�iu�\N<P�|���Ԕ��Un�@�1��iD��z����U"r,f)΅+}y��*dX������\A�D�� �Ù��ey�Y~s��֎��uP�nU��ʋ!<��L����O�"(
�D�g�&���ɗ�#��@�@�E?�����ᆠ���+@�z3
�,��E�7�+U�S�0�f�r�7��C���W���_3�y'R�3f�Q�x#�s������rWQ�;�?�F [=Ն��v��^֠�[�9�`���ј o�"GT�v��M����0�E�[��b��:��H�Xb#W�*��r,�7���m�zᙺ��~SS	ܷ������N�#k*�ж1����U!�9s���\K�
��2R^�_@��g�χ}�q�r����{ބ��`��c�R�6�Rj�]"����G�F=�e�]��W�PW�0�K'��"QM�1��M֎���?C��I'�U�'��w��[��b!]�4��M_��
���`����R�d�MG��I��۟�nm�I��9��F�d�Q��O�n�Fh<��c��@s������du�d�2Δ�E���=��U���,[��pvMf�o�=�?���~KK�s|�~]� ����kV�R!�ߧ��2�wTM'sv��m̪�(ӑ��p3�J|��VL&��S��0�)����n��[l"sp!���Q�zN�bW�S�sr�	%���R� ,�q��1n�k0�6���v1r�y��n!���d�G`��b��?�}nY��uú���2I�n���gD>�с3��7�1n1��,b��8T�l0\��k�v�y�@.��+nu�"!��[�w��9�jv�4�	�N����H�Wz����W�Vt�![��^d�-2r���L�����^�F��ѷ��M��5���h;m0vcO��h�D7OuHH��(�/L)+��A����O�9Kdb�*!�-R�އ_�
�ڙ���y�N�;��r���'�J8�ةju�aJ��K�W����=-e���"�Q��]Q�:�ɷt,1���/�=�c"�92�������i�Oc2F�ti*O{@7���K2�Dښ)X�6��@@�0�!�W:{p��d�
d#/��f~�;X��s�!,U���C�u�"d��Ȑ3�d$J͞<uy������P�ϒ�<j7F,YT3�����o%-���(������6G��1?٥V(&/~u[�l+�i[*(_\#7E��L	���{U6�Ô� �Hr��0�ْH���n����+@v��$!�C��M��"���:�[��L���?�&ǡ%����I����X��O�8z�'ogb$cfE���k���MV�@��yF�85�w�5�5
ύX���:U�gMjO�"��!�Z������$���]㒮��8�Y�x�+D�a���^�o�ŀ��H�u�A)w�o��}mw>Fw@�z^ϝ�R�M ����B�җ�gF����fѷ�?(A@/CQ��H�%=�by^r7S:T�)=����V����� �4Ck����aڬkC܀|�~ �$P�\-s�j��Q��l���C��@K$�ظj1�R#LA2�{�.�\u���4F��r#���L�{T៽|D�)ŷ��E�o�������u�m�F01OI�ʋ����Qr=�Ŵ>��ۊ��4&�ń(��CL���x�I�۩��h���晘�+� ��ǫ�&J���Y����ͤ�+�6�S��D��N�B�1n:���4�ѡ�x7ko>z��Eq	p�8�[jV�߾])_���r�Q��˯P��,�����22����R�s����7!k�X�Լ�����@r�x�'�2ٟ�����"[�4�,��IŎ�O� ?���O�'
��E���7�(e��nj�f��罽~���C����`YR���������ET�.cc�t@o�Ꙋ�ˬ�u!�\��Y�*������Մ��+��Ԑ��6�R��s����=�/ڏ��aO�W4W��W�:�F)/h��j/ �gi��!ҤK�E��Y.���_}1&��üh�n/4���3���Ȗ ��XI���hP�ě)�Df��~F�MX��F=��t��B��҇Z<	�1�_���fc��c��H���4d�D֡��)�%d���$��8ݣj��5r�ͤ�Ve��7��p���&,I7��'��h���7��BK�BR��pB�r�
�6�ʢ/n.2I쥒�_p���a���I��0&�L�p�05:Hv��0�Dռ�X�����%����-�-aU��͔�DZ�	{ps��B3�'� ����c��D�Q w��j�i��1���� �:�Cx��Yi#��p����]�I�H�b���N��W�~��Ӹ�o���	�R�|�������:@n���o6Ak��yZ �I8���@�xIdD+Kf��;<����7�=�bط�q_,7��
�	�zB�Krٓ����v亰����a�_)��46�h8����;H��(9��f�|����]��(>��NSz_�cF��P=���Nٵ��9 �]&&)�R�:�9�䙙�ME�����L��=�[~���*l7q����(�ōs3�1�O�N�U=���7�Dn�>(�ٜ(!*y�1�"G;���:\2[*Nsk0P�O��RZ���9iw#c�[�2�/�z.��"1�ӿ�;s�-ײ�7Yj��ٙ^���o�UF~ұ�c�g�ՠt��ܒ��M��,�f�����(�=��Z��^�Ku4�)�G�PMO�i�'6c�_�v,/�
� �$~�����sr��v��h<��x�r�e�����D\��_�`�W�aXJ6@���~{���b��>��˞(�榛g���4 6G6��,��,�|�R��� $KL�2b�x�pb�ti�QEk1Y}:6��p����)�F�{'!��ɭ�.�쿒R�y��;$�n׃���fc�]�^�#k�n��Vޯ�������x�4;Imv���&���7���*Y/u= ��N��G��q�����.���e�E����|݉�|$�7ş�Bfl������>	��7��:�^���8�x���#�O�dˏ�^��C�'ؾ�D�&;��hʻ=G�pY�������Tڊ��?.7m��f(j(��t]�؈��>8=�d�և�"�M���y����'���{(j0��[���T�#H�@��@o��u� � ��9	X9�>B��w�N�yrUb�����?��aZc�7�=3��ݞ�HC-�c�I���YOð"<�L��b�gnX��gm�
 s�4��od7��^Hs6=�hþ��`1?�P�JL��Ȭay�п��R[��ig�TH�f��f�1��B+�	~�'�A0�N0�+�����R'���[Se���~�V�z��.�yu�!��|�S(蓄��4�.�<�z����ߒO"G3?�}S���Ǝ�4��͐G�wLk���3�>����]|��3���-5�/��I��9dJ7��p�$�����\R��%���Z[����ʋ����<H�E�'N�2�x���Ѻ��Դ��B!�;��y{(A�T@��z?��b}t��^��Q�d�j(�ߤ����G�c���ܞK�8�s�|��ȁ	�����<�d�޴(	~`�2�lkS�>�K�͒|��^^#(Q�<O����1�� ���w��=�6Mn|W�d�l�u�~z��M:�;���#)��;ߢ�uD�Dd;`�u�P��+i>����K�����������W��pf �<(kthneΧ&����Ʌ[O�*V{U�������_�*��}�p7D/�0 T��c���4�8]`���q��������_�iJ��h'?��+yR7
�נmI�fR�nO}���ړ�ܹŰ㾋ʂ���(�yZ����#)S�s&��q[��܂�1h��}Fy�x���!r~��ԡ�2; 	��0��	�a��fS'G�~3�68��u֯��Qr�O"��
ʄ&[S+|����ם�+����;��?#����w[Mд���<y���;���j������\�B�=�A��;ʢ�G��: r]�3��)qP�B����ʮ��������1�;�>Jn^��/�n|�C��e.K�X��4�ů���i��H�5I�G����X��C}#|�M��;�ݎn�Q�4�h�qg=/�p`�|F�MW�g�rM�o�xݦ�V��ٖ�,=A_X�<�Mm���'�xBq�6�:&8kE�޷d10űܠҲ�*p�y_X���a$R���Cb�o�g/frD�)F	��p���'��׍��5cV����ц��z�Uv�'�]}ۜ:_IL��w���i0�gAoA���
C�HD�H���k��7ŒВ,�֠��d'���k��q�bF=Wخ����jlH��/�SY��3����"��*L ��M8L�q��8�'sm/%�S�|��<@38��m��t�1��o_ec���X�4ItuGQ�njrσX��l"�.�� �冨%��}oƪwG�=���!L���Ý���ZZ�	�CK��+��	��_K�0m�^���b����P&���vIn���kp��MK���eN�u��Mz~����8�� W�6�+��!Jn&�
T�]����>/��i�oc�z`V䄽�*���\�L�����k��F��/j��(���6��2�գWD���Fs�	j�=W��O��rg~W&F���;�m�������m��\$>[��L�ࣂF'}T]�r�����.:�3��a�����E9/�W�w2MY��(:8����>w�J�_#3Dn/�M�ݠ^��� z��e�V����Z�VO1S��s�RFYË����~��^a��&�!�f��6_�+�'W~��1t{���%v2���\h�+P��뢡�@syO�!���"����u
�}�:��z��LO�"��SI����E�{���7��|TQ=�S �����gZ��_B8�6��� ^7~8�I�Oim5�i7/�ۦzh��R�{�')�r �O@T���6N֤�W4o�%b�D;j���^��&#������@���kǇ��D# )�N�=,��O�Z-o��n���Q�"^vvs.����!f�$�: N��;�/*&��X��R�qJM�^���� r~jR��{83�g/³&x���q>J)�~���H���t���OjC��1׼2�����j�(X�M���"?�b�9R�q�#���EnY���X�Xs�<�14H�يЉ�J��p
��"(�N�����ayHp��,�ҵ�M���/�$z�p$uP���Sڬ*4Ar���~�{雰��� ��maa���މ���`��`P��4r�竞[��a��p�Zdz�{0��=���Y��2�S�V����B����,H&�e�8�@�=��Iy^đ4��ܴW_G��Q�V8KP��P�ѝ�0�$X�kݣ� ȝ�Y�����m��[�"�R��O�LHP�_c�Qo����K��@���i���k.ֹ�O�xߔ��^�]��0�myx�,x�,'�k^e�������S��x���f���2�5 �M[7)|"UU�r����x�*���h'_p	 ��3��q��O{T����fT+r��R��Chkv��J��:�1�Sg=�r&~C�D.	� ��&����O�m����y��+��ݒ��kI�75��>ւ-��4����5�C5W��z��HM��M�?W�/4F�,�^*�~oh�R�����<���u�m&���峻�S�N�Fa��j�s�a�� �ﶊ�B�h�H��G��Z�>s,�@!>fmC�Z=l�������4��Ɉ�b�-�I ��7��(�d�w ����n�N�K�٫Ts"X��$�tc ,�yE��W�Y:nBy�ak�m��@��K�W0e�՘�ЙB�ͺ�Y�7<s���,�n�gOU�d����?dk���,kKIr�T�K$^��������rNQ��>9�9�#3�q���a7C�����?
=�~MJ\k�� ��.�H 2��C�W�)������(
���f	H�����2��.�G�N�ä�F�'q�� 7��+TE��fL�Ix�^8���]�Dr���*�y*jO]�8L֙���؍(��bpk3g�wc
-�G��S�wK�oj��(��Q͒����o��}D�D�3�]�_���,���H�V����ڑ�{ז�����?��9ǆ���M&n����q�L抂����E�@�ĻZT�Q���݆�__�c�mI�l[M]J��W���&�K9i*̺��/ME$O�&N�S��eb�a�L���|C+��K(p����PO7x�e�o7L}j�L����bY�Oݐ�<�?*�"|8)?�`�6C��V^(f� UM�A7���#�H<#��T��\�-����ѹ��Ak�;��WA�h+�#�aiօYo�j���O�+�
WVw	+��{���@ �.����[+�ֲ��L��ym�b~@`E�kBh[��X��&s3ūچ:=M_
>�a�q3�������B� �
?�SuJ��fگ�Vې�g�x�6���5��:�DRh̫��x&����p|����T��'�����i������<�5��B��i?��@u�)di�#D����@�b��؆�y�ڝ�,���8b��z�2Q�\�8}wa�rw1��m��j��o��\@�{�I�V���Ӏ�k��p�D'�d(0�.���h���zN 9(+�-(<T�}��.
��!Bj����)ĵ�z`
u6���c��eLIQ˞˄��iw��L��c9)�T�x7��h�;�m/��^b����~�zK���`�ԣB��I�^���F4�i\��9�>���;Û5@�s��'&��f�
Vg����l�Ch��6�v@�>_-�_��0K�M��e	��0�J�ݮ�M�G�<^�0�m�H�@#H7zQ��Ra.�{�V[���F�7n���1k��n�[���R���a�c�mZ�~܄3\MYH23����־~X^��+[d�o2����!���'y�`��B��`�H�HGPbB���.zQעk
?����o��� ����P^�%�჆R:�%��w2�iYRK	FtF��(�I�	~�	 '��:�Iz}t���:;F^��*��q����æ B���C��ef�:L�HƗ����,�#!.q:����3�ʞ���Q1�(�B��0�e4�$��6������1R�xsT���@E��}�Y�5O�	O��*
޴q^�2ڡ|�0^="�'�@�~��b	z�H�5ogد��o�{vT�}��t��)A�и<�|��0�+�-�-�1^;�7����1xu
τ�=Rꎦ��O`�SHl{���0�Cw�a��eG��+k~�D_�F���Y�X؈|a�y"�%1�R{O=���U�Ҍ��� ?�_H��{�T3��;M:��;\�ʗ������GA;��c�Q��m).�[����I��A_�{:���<�7�}2VaR�}p��8yJ7���)�v�<x߭��|l��� )Z��5��R��tN�u�%.*p��Powo閂Ә[&f8��҇���=@6/��s>D�l���Z����.�y�:5R�Cqΰ� |k���ݴ�=Z�b�^|�yZ[�ˀ6q&O����-#�!ɯbf��"L��Py�h��O~�Ou�3qD�v��p�9R�dg(j��&���em<�����3��?��Z8���tHn!R4�'��Dt�������$�_��|>)0�.�P�$\H�TH�խС�s&s{�%�����1͈}H��dyL��t�ſ�vv��s@����W��U��P�MB�<�<���	�r�2��n����|{v���S��۳b>0{&z*��FW6N~A�LK��N[�<�p�Ѧ��P�����K�U�a�Ѵ�:a���� v�����-B,&��e��_����,�{˴��r|�!�v��ıX���G+.F������X�*A���phcM��d��m¹o:�%�2ȑ&���{�c������T�Lt�m����ݑ�@�o�W���W\T]�I� ��O�5Uz"��Q��[���MU&�GQaײ�[�:�I�V�Oe8U8D~idl����=]��ՎJd�R�@��j��2$-��"q[��^��k4�O]��]�0ֱތ����4�R6ci��j�l������V�P��

�O�U�@�r5Mm�7��I��3}��i���R���X.�?�ŋ���~�/>��`<�\�W�9d�"ݬj�9�� ]����-���Q�B�j��r܇B#@6/c}���Ӹ��dk*�xaB<�-5*ICR�UX�|L�̯�-w���Q�wA�MO��э����U\���)��\yӾ��Zģ�gv�c ;�@�-�7�1��R� �z�JK�@�^�m���:�Hi`�TYL4}�Fs��$㻼|զ7��ҝ\TC�$�Ł8v!(�paS������g$�fnq�A��\����c1p	���4���=tQ|� �7���	�����[�*Sůˁ���j�u�e��v�Oy~�D��f8d~�>k+�$-V���ӹdH�o9�/!o�{��,���!�[C�V���i*���(�a!�'B�IR�]���%�o`�[�]_��`K[N�0��7l��S�B =$/�g��۔	�c�胼SĮ���/Z�)7K�́���7)Q��j��	��L�m�4r�cT�Xy�t�f0��c�fq'� `V|�5��󳡋9v����lޮl
����+�gM��a�4,�n� �����󺯂�AP��t}X���ˏOW��ݒ�FXl\��� ����G��.��u� A��`b�%~�Y�9B��_|!�i���"�s���p3�1���KWD�D����:Q���?O��aD��J7��0j�"��3b�`��7hP3��Y�{,3^1�a�k��R'�7�Os,=�Q��=�,��B�:XT#3M�B]��3�1V�e1�&�u��t����k�U �x6n��yg��R�� �<���L�@�9d���Xl�73R��3N��~k���<���c�tJ[�/�� �k�T^F�v�CC��
[.I\V>��P��ԝ�uWqQ�1,�b�Ҏ8�=�F�6� �w:!�W����d X�L_�K�wbh
��;ur�!v6p�Р59)k@�k�co���V0��;p�l�q��t<w�� �g)f�UYҢLo^ ҵB�mX�5�Xa��H7t���%V�&]��S�b�3⽲wuD_Q�؅4M#K+�E�b�����Ў[dH/�X%���=9��L�,ט<s��ٮ�6̹+<'v/�F��_�)�|��	7�ڷ�y���3Z�nl���QV�8h
��8vv U�J�E)ji3�x����T_�z�K;>�1E�����P��r�FI����#@�}Ί�I�O�>+�X�n-Y�G%P�?e)˘k_}U$.|O�xs��x�@l�O�Q~��hPI�u\�5�-N�P��aS�{}�b�\��:�� �D�{秶���訫Gm44r�AOߋ�|��Nm�,��ZV�A���B��Ǜ�^O��E�#>n�i�g���8zǚ(h����fY	���v����Y�:�'6���|�giّ%���H��9�N0s)ќ�Y�g��g�L����3��9h��Q+�������r�٣��J�R:�/2��[���4�0z��V��4(W4� v̓�LK���8e�Ig��E�+���7�`OY�G��gtl�M\L�g�c�����μa�0�d��2C4$�&����{��	g��3'@�~�d/� ��e����G�S�Pd��#����
,!ϖ�g�����4�}�{Wՠ���&��o߶�sҦ�%O� �g����D#Q�r@�UZ��lg�o���]����V��ma*�6���҅�N��V��\��������#[ڲ�D�nʝ�s�# ����O%�E����͵m�-�`����V�V;���~K�C� ����xon�F�X|���B`pkv �Z�b�8�܂0�a�"�ć���z�EXE��� ��*J0��Ig(���v�9v���=�g�!&Z���	��pc�Si���K�ƌ�c�P��H]���&��@�(%�/�#��%�Zl�/�5k/�G�����X��Sh>\V���'�p4"��9ud8+s_N8g������� r��ԡ��(�T��[�����I�<<�(��Y���6(2D��!#`H��|�w3���F��S�ӿ�ǒ�*�u@D�D�]�°��O��^�X>X������{Ī��P�,��tY��W�Z,'F8��
�B@�sKXy�gɜ���/� IA#B*k��%j�JC���~0���]������]U�4L�c�I*}�������������u�%-�=��X�LM�����z�~]�L1�p� ����EK���t�}h������z���ٳ���"9�%�`�mT}��*�	G$��1Y��~�#�J� ��SC�ظX���s����rC�<c�������$���;7\w2�� ��߫�	��L�4]W�B�L��m��>�U7�<% �c�z�Йy�{EC&��F+Tq�m|�?/����pJ^b+d/��i�؁[�E��YG�����ߎ�� � +PG3'�B_����!��&߁�#Jh��� �;;����� �����/}���|Jݦw9�.�;�iw���M�9�L��F�c�o��r�L�#���1?L��d��_�i�h*݇�#�`�ح�7Q>1��B��ǂ�L�LOդvo1���t.t�7P��1�X�-��%!b��>�V����0�,�X$���	�*֞�e.TWO�x�kaB]���O�Gzb� ��0��l����L�uP��\�ǜ���E���x<<��pRc�x[+t�g�C�`�ϰa���bf�&ӈ�?�����s�U^� ���b��,�|�ނˈ.��R���Ž�^��Z�㾡�����},�@������"8_%��-�����-�]�+^I^��M(�_��{�?)x�z}��e~��4Q��>ڿ8�/�j����!ܙ�|���B��q�@�|��)�7��H�u���W�nG���{M���QVȖ�8e5A�Zl�8o|�_��8���:�� g�yI��PBx��/�7`˱d����3��Gp��S��!�%�Es�K�&�M�#��'�j�/N��<�Ҳ�1��Z�j_VI�j���r@��,����&�J`�Yb�<F52"����Ansل�b���(z�x6%7�S"	넴H蹥��J\TcJ�Z-@��÷
9�Ԣ#��3�acWR�0��_��5x8\���� ��MZ_z�8
˛^;�?֤!lZ\?|S�WL ����ζ?����&�H�����1&=f�,�˻���x��T��KB�&��u3~�w��\HCM7S�H���^��)'ϓԞZq�h��wr��x�nⅢ9u狃�̀�B���њ���k`�"�����~�́���i̼�B,�ewM�%nZ��;��k=A8��Z[��o�\m���}�/ E��&��*=Q4aq�;+����ۡ�.:�5��?��4P�uoQ��|�SG�fE�6����eĥ�xDb��|�ݭC9�k� �ə�����?QtD��ENVL0���N��~�+	9:��+?�Mh"���"���Ia�E��}j�O��7}$�?u�h����`�O����-���Q)3	��"���<������Sg���͎_Y+���*�_K��[�G�ˋ�vG�@0b6�cR (.������̿�'>�=�clҨ���hQw���]ܴN��E�&l_v`����4kA��H� �[,|q�{4�b��-%���Yv����"� �]��Mj|�;�4�~��
G����27e^�>0ށ-o���~��+ssz�FPj�lD�y����K���)�G£�u�ƥ�4[�	߹�I�Y�:��d傦���C�7d�G�W�ep�"%�����7��>\P���N���˗�-�S�U��F�=y�UR�Q��l��1��9%�C��Ţer���2��뚛,�ί��/w0�ҙ;����̫<��eB�W��P n"H��{T�E̳�1���ռ,�� �Gw����ST�w��z�nH�<5�M��%�|�|3(�K�|�,ZB�2��	B���EYf�FpV���T���0�9|vs�/=����ZN��{���!�������xl+���D-�6 �7M��A����&ӫ�`�����1�:�����f�3��u��)j4�}Ss)�M��R��nª�O�����n��=�.�D��e��Ɯ���*�Z�
��٢���r~ ����_;��j&oȚؑ��wȴ[F��J�~�Z>�;䂛;=��}y���*�;߶�wL�����=������U����[_��.(�`�Z�Th�ՠGg��_��KZ�'��9�8l	N��Ѧ���в7$�C�>�S�S GhBv[�^��ASo���tn�7#���Ku��@Jd����r ׶s��nb0~sè���X�D\���x+?�3�#����n�9���o�������a�w��*`5��B��9�>�H���3*�F�����xX��������2��3��� G� 
�t~�e����K� �l�a�JF"4�]e*[@���~���h�6W�V�`�c�U���)D�B�0�]�k&⨦ �Cn�����tewz)�s��3D7�n�5-NϺ!e1�HL �a���7���Q���S�\Y[��e}P�7���i��2H!�Շ���Hct�ʌ����da`�3���7@ -�F��N,V
�p�d�w�Z����kJ2���Ǆ1�M���n�]%[,p���~���ظپ�ւ7F��H馀����F�v;�ې-�
N.3�V�eh;ے�	�/��/��1�M�Gv3q� �JB��$	0����wz�r�-�n��w�P"��vw���|��=��2�:^y32E0!q
��ޯ9CQO8,��g�ǽ�@$��p{Zo�(�$�b��H�oY����Cd��� ��m���1�'53�Ks��o3@Q�#����n��}��K�;�������'�1�T�e��$�lo���]9M|���f ����40��v��	�?��f:��dh��|��q/����ɗkցF���1o��%Nb���h��#n1�Nڲ���BHH��%ж��/�9�2����?[Ζ�n3)=��LD0sۋ�8��������������f|���4ԛ�	�?�o6s����;*\F��gE��G���:����U��r�"����3��I�*�*�y-�~:�b��=�SF����	��-y�������8�z/��IzGq����@;���AT<zOJ���ō �{S`� A.��A V>B9�xIF}��V)�C5KaPa�o�l�Z��=(�A��.W+�����ӳ%j*�́>��(���O�������2a%.�#G�1�y����ݶ�&���K��:�d�]W?�:8����h`����5`���q�#U�OPρ;�P���!�aԗ2S�]���1�E�C�\q��z��oN�K%���OEQ6�����F���&G����<�fx(���W�;a2�����`�a~:��W?�i��^�[��+l�FgfhĪ��ϑX�rO��w�1�kկ�ܷM!�HIY3[̶/�B���0$�� V��Y@��������Ǧ�Qpl��ђ[9D6���[e��Q��t�'�Wyj��XA�q�Bz˵�j��g�C�e��(-CR�����P���C�����64�)�D5��CGY����X��ˎ�nyg�p�~����7};V̀�+�f����9��%�1��^�$�����Ɵ;B}�Q�V�3�*4C��&NѤ�0`ڧ��˹n0��P��CW�"�jL�Q��M}ZL�h.�<0�����0Z`�A+&>��Ǡj�;?���3R��`6�����\[�!YJ�p�.w\z/��q���E&څr������VGʓg*�ّ���*�w\�u;���Rߵ���l���}��A;�OF?f�xQL"C\�;(���e<��u��ć�A�����@��D�"�ن�۵�����WE:��^�l�׬}���r������h�u���&��oټd,������b���)!��"*&VJ3(��Q�`Y��S��Za�Z��+3��g)�q;�u.��I�:KbC�&�**=��N���Aj �I��H�x�w3����e��L��n�=G��ז������2�+�����=����*:+��̄�d�U��9�q��'6�#e8�gᣘ"'-(��-e���m��[�
Rz:�0�6ة����&2��sN8k��{�|B�\�,G�'��x��'ſ��Ml,0����V{g�~���p~5I�A޴3�Bȩ%���"Z[���@��A���&�R���-�t&Xʔ�G<�Ҩ �72h�+z6�\���+a`��"�|�V�*A9m);���,����h�!(�	 "޸�'�䂧�R�	[ ���ۡ��:W�R?�v�췪�ů��cy�җ�?Be_��:����]�g4 Ϲ�ه�n����
��HE4�n�������L��|:���2�����h�M�j8B��p�E��V�d���	���
�} �P��u����������~�X��<Z�H!��)�&��ެw.glR¢}�r_�P��i�>�Gz�,Y�
;�׀��A�����@�H��m�@�f	ŀ�}d6��r}��#��\���Q妫G��BY�\�����s�\l�����ܲX�R������ OZBӁt�R���i�M�>�-�躝����J�i<Hp�1,���ھ6DJ�@m'?;&yڣNdw�#��z��^Zh�h��P2-��+��+)���BB��v�	�n��4N��^��ӵ4�ژ�?�6M�͑n���Z���W?`M��W'�mK���q����$�Q�Kg�/�RF�*������SD�}�2�*L�����i�k�_�#�����,������u�p):��bSc1S�A�_h�hռv� �4>-��4ah}�wި|��[���E� �`���RL�k ���5���%��x$���>�zL1Â���l��"4g�Y��'L���y;��{\8K�[�"�^��P=c����NIH�}x�%�c�c�\YP��6�c��;���S;ڠT�@_ �]���U@.��%�����/�"=�4Do�r1�=q�h��4�|��_B莶;�o��?)��#�^|�Γ�r�S̍yoG�(�B�^xB�z�a|���4�c� Y6���_�����T.�_��D��L{d�N�eU��z2��.5���m<��wy�W�|W��,<��5����fր�2/{?Xt��-�VӅ"�1 hy0���?F弆y|�Kﮣ�Fb��C�vA�T*��I��l8�Lݍ�:&�	��ɻowC8nVf��rh����F$8k6�jlo���L�k(�C�b(��ڬ%��?Ŭ�Ʋ.#���N�_����)��R{|]S�3�ܓ��6��2`�3ǎ�$yO��m�ҷLA&n���?�붸�4Ҁ3��b�,�7����1�E_kX��uF��)oTX��Ȝ4<1`G+W|:��s�{<�Q.<�%C&�|���i��y ^{c�><�rZ�C$�}��{H��q�L��0A�@�cE��U*,^��V=.fäS� _��I�P��I�z!�uˮUz!���c������,��E��^epׅ���n�m,Ⱦ*��|�DB��s����G�<�Y�F�k�r)�ekam<���Y����K[p:H�.Gt�	�	3I3A�ߠ<�9XRo�@�{��_��bWY�U)��U�d]��i6W6� S'�oJp#m�Y7}>H�C�����jw�l�|ۡ؆B� "H�Le��]�xW�u)+w�D�~a��,H.�Z
;%�3���#0���K\��Rp>
%u��0QY;�Y��ܸ��//�`a���2���-e�:0N�0�]J�vZ�3uEA���_,z�@���0h$��IfE|��8��?i� I��h$�"�'��o"����������q�{p�m�b ���>�y$c&�݂E����i
�[��`	�sU/&��Z�a�%�"���I?�5�s�w�۵����q�vFt���y�Z�c�z�j����j@wX��2�5����1�T�D��'%H������c��QW�A���k���H+#�����Am�4)?��$	�{`pD��*��6� ��	���M�T�ƽ߾̅}���=�c^�1��T��������������y�>e�����cu���.*LM��k���*�]N�����'��D�k�I�*y��VK�1k,��TW<\�� !�*�_R>F�6�jȖIx�Ϣ$h��`���P7�#��}�_��_�\�t�`����,HL�w�=
G��m������mj�T���<��h�2��"��.����'�Wm��K��,֍�p*���&�_��"ݾΌ\�����-3ߧ�	�� ;$�"���+��&�Nz۩��U7d���߳�༱l��C��Xm��{' ^����r�W�/��(f*�+�3ߴǮ��R��1/ʚ ���8�93�x	|��hO�����oN1���fO��%$���؀�#w]p}��߄g�h5.D��}�mԓ=_�<�y��6�~���}����8yH��Kq[7	"ʆ��(&��B�E$$Ԁ�ȇ��z�������!��7�������f���.�.It�I>�3��X�Wv.�\(� ��&L/��+�͒�%��>�M��M!m!c��*�8l�/���m�b�TGofj�WH�:��/���%F�V��8�ˌ�1.7�cvh��P�y�N#m��U��	O�\�V�eh�V����u�(��� t���}�v�Ρ�[2��v��%_\ �w��+���2�`�r��d�S�|�H|Y0:��}�W��'�L&�i�w�ʯ�3U@�-�RV�ʉ1�_.1[hvH�_-��� g�JQ���ո{�>�X�t�* ��ޓ3��W+@9꼡����ҫ�	ba.��daA���TY����f�:�~��tZɜ������܀�UAZ��o���X�	>�'&D��[|U�.=�NQ����M�ev\�8�+ǚM��;�}6]Db�$�p�Vbj@�!U����H&�ČQ����ҫm����7�
6HD����Lz���B��g�ݼ�[6UzK��Z�Ă�Љ͂�d�3,���m�"�+�xP|����1�EP��N�)p���KqPQ<���Q�ܙ�����!�#����wl
"jۡ�6��*�Q]�^��XWo	%��~�<���SEED�Cʵv�H��R������ �ɣ�����P��>_pw=�CI{��s�c��i/�/
Q��O�(!�a^�'��kD�P+u��z�:��Mj�Y�H�h섇����/�*D��3�5�-lN)J$��X2�;O֑'6�)��ܮ�� 4��I:��n��[DP�u��M\K5����=�ڟ����_6���+�~޹��<�S�(����pU��i\n�8Z
�� ���s��� 絚�d�w��E��,��徠���f�e�;��]б̌'Q-�j��&���4�$���2���S������Y�$���­��`�XY�9�������)��q��6�omV��#��R���{B��������x#��q���e��6�
��#Ƽw�4{�[q�����*�����)�~���e���ZH�G#o�.�I��V�V�[���p��Wa�Y�ϑci���9FϜ�{B@�LO��;kX|d3E� �}H���9AX���GBg��$;h����= ���7a���m�37u��ë��e�����!u�QXc���	+)�y'|]Y[�|�`�c�F�$��Z�k�
�kBl[|�"#���~'��I@X�R��mX���32��5��K&#�q��ʹ�+且N_NՐ��b*��ұ����4[q�^1�n4!�"莔�Lk����i���U�JCÀ��SX7x��%zZ){���0D�XQ=�\�_j���u7G�>��iThviX����xE߲i�[�����J	o����0ە��L]��l���� ��Wpa|�	��t�����iHZ�L~,��8��1;��ȁ�ӗ�N��<u8F&�x�I�d���� �3��80n'p%*���v��hl���_׌щ��^-�8n����BO�t�C��a���C�͜0�3 }��h����c3��t5i?�qye���T���Q�Q�KT��.��#��hO����0���}�K�;�⸥�p��������ª^f�UM"�r�PE�'Ra��|���'�������:��}>NMGO�����dϨ��Ky��A�dD����a�.F�J��[⇂�L�#��H�dK�_`m�2��*;�w݋�
��d��Sy�9����d���G'#
5�T�n�|�Ϸ�~q@���A~:ȫ<k�h'/#�Y���9М'���+�%�G���W��''�� %�����m~LL�ݐ�ȣ��r9<"$0�����1��XVLש×>��N�.j݇��2��K�c��˫ʶo�� [���&0j
��s�y��I����xb����k�X%�~i���,�SQ�����>mg�IZU��݈ڿ�5�cgò��s���ON�G�f����غУ�LQ�ԇ��[�EL�2������I`���n��@S�]dd �_/��\2���~I���Ч���Ѽ�^�X���:�-��~P`L*���c�9���+w�r�Ҽx�Eq<��l�A<����L)���uRb��AVN���`���l��nv��p����H���q�Y��v�xv��yf��GF��ۇl�N��%O.��*�.v�g�_�҅�c�pN���F���Օ�A��^��
I��+q�]�h�M�
�4��yf���u����FI����q�l=�i�W���W0`MC��%u#�m���|�:�[¢ňlA{T�N��x�#�'����ˮ>ҁ��.�p�� �y�iA��Yn��w�;�{G�H��zk-;��p�[����N�]D�V#*����'��H�����_E�m�K�o�� x���4��o�"=-�1�Y���'9:Q���n�Y/IW/<O�y]2�H�5�����i�4c�zbpn��ՖM��""��V�+��U�;G�aA9�}xbEzw�/��k ��]�[N�}�儌z�I+I�$9l���xb�MP<�+�?G����6�&���y�08�~�������5P5�E#'Ѷ~��3���/�4����U�g���I5i7��%O�o)�(�|F���Xg�~���g����|��:N�ܢ?k��D�C"2�����������]��x{�e�>���X��-��P���ny��δ��<R��h�]n`ZB`��S5|�A�m1AⰝ�@�'�����!�j*&��x����;�Ȃ�iM��?�a �ۚ�j�x�8 ���Xa��bu�WS�g����S���֣�]wZۯ@�(uD��^�qVR�.9Q�u~���+�d=����W�vn�|����@I��|:P-��1x�e=h�8��꾎^C��l��c���%���H`{Q�z:���p�d��=���{�3���K�""���Mw�������)(0��)�|$,{�:W�*�b��NShݘ���^�'��p"=7h��{�ӆ�E�K7-4��D�L[� =�XJ3���+L�D:(�v�������;ˮy|拫u�%i+G9�Pu<�G;��D��e�F!tB��%�[�.�5�|ĭ"�!�>������yp)�-��FT����vDIz��e�{���3�(�%�|�}[qotĤ(Ϲq��
u��4&���+�-��}2D������al��e@�?,7�@ql���Qu�YD'�Pt��K��#7�b�; ��+��b�"��b��
!�[eV�#a��Cv;�Ǭ�0�"죏� �]A�^�Ց�i����6�#I�j�{Z`i�ɱ�^��d�<���K��_��E	M���2U�Iܲ2�=��o�l���@/�]ˠ�yt0>�ɾ�� A2�H��zڠ��+=>!��S��T�������p�E7�sN��z�Z��?mOq)���N�#b��g.eҘ���6K^2�]�����.�s�@�t�t�ot$�{���8B�t��br\���D'���k���BQ��#[��wy����mY�glgj�(�'RA�6��
4C�!�2�e�M&�P���n]���詼W�6c��p��IS����"�GU�x�	#y^��$�;_�G�|5��vx��oW��B�z�s9���. =#��M�0������Ho�����]��_)��J8���^S�w���	%�jK�$�L�qB�8��,Q�/۹%l�l�x�c���B��0��o@еiH�d�J���Y7�uI(���P��o 8��O�}3a������ᴑX��P���a}��a2��4�Ƴ�ww�}��p�bc�&~��a�L#�8�+Xh�zs�â� ��@��<tL��缃J:��@wZM��T�"4��ȤnT(�a�=G����� �W��x���P�����`B{%Q%R�t��X������T=Zܴ���>��}���3����mJ�#]T�����o���,�_���,b�C�"�^e�������^2',��5���bPwy������vM����־�>Z�����Pc�	��d�¨����%�z�"$_>Ԟ�������5�T���(v/�.�Lk�	e�&\���x��zs���&�ǘ3��¤t�q�1Գ��*ooE��+��`�v�&8�aV��O�R�K+Ih�R����" ���	 ��^"�4(�w�(��r �eb�%�A����f���%`"��wL����=%l2��C�R�BW�6F�k8�]�5] ܚ~��+XY]��AK`�����PM�9�~�Y(��qsw���ڄ_@u�d��f���PO��J�����Q?hΪˎ/� ��Q����Y�i^<��W��/�Nыbct˷ӄ��6��iC�
�W< �0�~U��wU**
�D$~��z�J�!��;���]�2�I<H�D��[c�� �v��E5?N�>�����_b���j�Ʈ�^�9��ie>�����+Rjշ
�!tw�=����A��}�EC�J��TQ���O�ܛ_��M�T�۰�{7vY���b��)�@�38#J��'�~s��*B}�Y��G��MI{>��b�|Bʆ��l��nM���^ h�,�B���o���4��m�� �wV��,�Kϡ�<T���_��X�d�?P��i�����`�*��Z*r/��-���c���3����Q�C���d;Ы��b��ה%%Z�	A:��Ҍ�ta��YQ|?��*9�1�G5��<�Ft;�
!4)�X2�,Q[0���1��h\�v���c�Uߘ�?�o# _��^�0KTgy_�@�"w\ۯ�]����C����&���aJ��y�/�N��m�/Tb)P�)��#�O��^���2��0k�*'��n��Z Y���\�������ZЮC�F��g�j�ΗJC{iu&R��/�w�F��R�����5�g�pkZ��~zGU6\=���h��:��H}����؎P��ZJ���5r�\�g��� vDWmW��iͯ�x�ڴ��BG�W���+�됝^H��#�.
�;�/'Ժ29�|6�M�^�X���.��Bj\o-c)�j�x�3Vk/X��L���0r����ʄ�����bB��p"=�0<;}�~B��k1������'�b�I�*��_{�h�e�q��P,Ҭ�e�|zU�#��Ra�W�گ<GȜ��t���t�z�e���f���S�`����2��$PCٸ�	�l=P������i���et�8g�����ď�e�I����R.s>�P6��6��z7�c��,z��)r�Go�%Ȕ�ϛ�07����~y�Fr��[Ȥ��؞WZ?�v%o����¥-��^�V�k:s1`�s�~�q3�9�bĩ+��`�N�Lw�P�2

J%�kUz���#�~�'����-l��j�ef����i|����H�3�^�= �}�Gc;�&�����'>��fD{O��f����ˡ�⡉��z]x����1���xχg�5�t���V�7x�x]�O�����KҀF\`.T�Z�RK����D'��9:��X�rI��g�lXD��uM�GN��$g�>��-)(�%��!Xgv��ow���@���ޟ7�92����D�gF�U�}b\�(?��*.�,���Z}�1%�9�m��v��0#�<s+��q�rm�-I��	#)-���}�Ii Q�����̛��,�
���1�m��>Z��>M �8m̝<ޝZ �"��J��$���'!�����>w�ok��!\}?@�vJ�pI�678%T��"�N;0e�8��lnؕ���:($-���N\E���6�~�vZ��R4�B+B�P��"�a6 �[�)��X��&��b4A���)�(���ʤ��(��U�Gϻh��#����;��h�j�+ >h�\�&��G>v��^l/ ��N4 ~^a����¥��OxFt$uٴ���'�.�d�@Hn���(�hי~���>e|�XW��
Ŝ˘( ��df'�ܯ6g{��gh�
��������һ�y�`r$$1_����W�Z�Jl0�	�y���w��ф�%M!����p��)�˲���9���J���N�Xd�K{ݥ���F�h�N��hG�Y���m��E5"j�oM�=kh����3����-�=f�[Ŗx'�c{��^�X��/����7vN%����4J��<��l��_X3�F�2�y&k(�;f	� fy^�4��l��j�~�8�)�������F�@�Q���Vז���k5Of�H�)	��eU1���#�L����g4 ���&>���=rԻ8Ԭ�6mι>�w��+9�x���b�ֆ�71�.Ɇn��VU�3S��؛ݐ+����(��8��ҵ�zҢ8��ʞрB����?as� _��:���W=xN�~Qg��O|��܉��"/�]����g�ZpR_�9�e��5�������>��.��Pw�#��\kd��G$��h��]�֩*.T G�"od=J<��4����֊|w��hj��-NL����R:�Sj�;Zh.�V|�2�Y�?W��yr�z�
��Ùj%VO�u��_�������D�Ǐ�� F�"����{]�{K����6���z�}4�+���q���9;B��v��o6�������աчzV��Q�0�B�In�kQ��>4����D���α���&�>����T򬰓�C#��Mݖ���-0�._�m��z%�Q�g�$wL=;�rmU	���WSH��\��?Su�!��	��/��!UL5����7�=QQ�ÊѴ�]�'�Y�I�Ck��-G@p���"��9#s��Z٦��i3H��jH�L�5���uE��>��Z�����؝�"�K�U���v�/��R?`���"�ۼ:�n�Ǥ�W4�w�܋�YU�wí���G�x�')��qN��"��k3݋�%մ�(oL�����E]��/"n` �ٸFJ�g*�(��IE�͕P{�x?7���r�w����0��T��~t�S����,l���d�Q�v�C�g+ff��r�b�H!�Q)I�E^͑p��5�`?^�����?��i�E`�0�Tʰ��j|7�q�����z�-,ɩ�iV9�D�12"=��xk|��z�|G5������5F2&�4�v�3=z���)�.�%��
�h͇B*%����=�E�f+11��(7-��~����t��P�!|��M���>G��Y7��[s��G?�~��z}���ޖ�j?���@�f�����+ܜ��&Z����)	��7��v�A2A!���N��*?щy��$%_�bs=�Q0����	PZ�љ�\�ωf>�c�z�Xڿ��%0���=��11B=�D	@<��EErʑ��x#��>^ըe��1n캿��A��qeƯL����6�h����Р�av��\ގ� �橗���f/�����4� �4�#�,
��vX�����]� r��
��:�׳�i�����5~+	u�t�$y���ԛ<�)�j�d�ە��<-U� ˲E0��U�,�Oʓ47~���A�I��wW-L��
,+W`�}�\@宓�X��T���^���L���2��/�Wc��π�)�5=s��4
����p�~�\+���L����j-�G�
pR$k��c`e�W�剦��t&]��H��<4��>�QVs��:�!�����Ny��U�U��|���$���'+�N3ȞH�kW�fT]�����uEL�%��,l������0u��lWN�E,�cHg�EO�M
������CQ��tE�y�lf�=z�'MYO�n��jh�e=ul�E��WĆ,��⚟�H4^�%	9�*���F/nn���NS�����u������_Ӷ`�Bhm������ޯ[$����#(�i&'�����wT�*v�4��nc�H�}u"(#c��9Xa�l��UZd�d�"F�S߷bBM���u�������$�5L7F��W�f��Kv�=��ލRTl��h@���6O/�8��c��+������a3FK_��"^����JVbJ���g�����igѢ�lֹ-��AFJ��_�Uwy�@nVj@:5�,��kD1B��8�ʐ�7���	�fW!$����������;��B.�]�d3���]�K���jvP��9���}e�v42�`	L� T1D��]�+憘O�b,����#�9e��Q6M��T%�x�yE����N`����j;�:��K�BQ��^�
��;���P�Xo��;����G�}("�a���lZ�VW��< ��>*�ȕ��:�V��e9r`�G P���XXUv���;�jX&�/��9�͒�M���C�^� �\o�`�<����>��w��6�wb� #bm�]Y�&�d7�ڰu�۹�̳5�2��t��0���t�Z�w��!�*���њ�L�:g��.�E��'��ޗ�FO- g���f.S��-Q���M��P�@��⤶���x�x{2�yN�y�@L��?�]j��f��ya�9�|pj��BF�CI��K��-���[S�r{d�x�cA0(���j�=h��e�WA9L��^�(�v���rBoV$��&�A?X}�g�W��8�J�
n��(Bx�<�G#��
U(>b���d|�g<�p��Ȩ���ϤEK����$i2�%8 S�% Nnol�l��ƕ$��1H�a��G�|PN%�|�u3��'�7,����x{m�]�'ǟ�>���l�ΐZ���S֭	Cuх=ߠgeO�}���G%1�0�һ���!�� V(�7]����$G���bm��E֍��w�paƐM��y�]{v�c�МR��yjH�P)�M���_���f<XȌ����$HW�)<} ��Q)��ꀥ�ڢh�ݬ�:r�v�f�`����,6AS3�� ]�j/ϒm�*"��,������<��c$���S	GZ�@D�s�6�v2�_������`�q��z�|�L��*L� ��4k8�&R�F̔�Rj��
��=� {Z���6�����8-��.dF��'t�5<5#�-��U��*q%���!�?��@�D��Ui"s����F���%�ڲ��\�|�-pJ��A'ϵA�J�
�$��*W2�o�&儲�������6N��C1���6��/�%F��.-���S]�q�/o��`d9�<�S�Y:)�|�ڙ�UG,G��D�G���H ʤ%a�'���|��&�����&.�n�� ?FF껠/���R
�(�G&ڙ���\�	\�P��������_�<1,!V�H�#{+�"\*�� .�*�Q�M��"��az�w�ưj@j�ם{�Ҿ<�FK鱬/W��[R�2'mP��۲T�2t��;��j9:'�8'�����C���	�xN���p�KdL�r�*�*�19�8#�`%��1��%㝏�R{�$��K��>K�/p��3���R;�t8 ������Κ�b����D�˝��� H�H�u��8��D;s��k;nظ(�|:^�&�J��P�wi���'&����R��Ա�پi��d�c�yƲ~��V��-�q�[����1N0	�
�u���/�m�9*���FDe	��-�)�b99{VH������:i�Ozy�S����݂���뼻/��^t�O�2�ɔ��Vv���D7��X b�]U!��#���<�������v�>�����Ĭ!�_��}f��A̠�.��Dш��4�S�j����m�`��p�'��WQc�c���X$�քY�������oZO"+n���!s�ǻ��I���%�*��X�Y����x��/�� ����"��kE�������C�l&�8��TF�ղ��j�G��KãE�p����£Z�����Ț(�łz�������������<����I6@=`D(�~Bh먉zA'9�u0�dc�mQ��8�l��=�E�w�UK";�|&ڗo<ga�D�ݢZ�Z���ȟ�+�@5Y�`��j���t�wL�洪����;���M�4|Aް�'5�+��¡����kio�8��U�3
�B�S��%�k��Y'a�C�<!A1��K-�d\�J �Рne!>�I�9]�ِ�f� <�SA+���e��6�S�jy侌��
 ��wOYnc}]�W���@��x:�C�g)V2/���ݤ�ϐI�|�L��޾~O`U�JC�L���H�#�
_G1V���gl*�|ğ��Z�b��6��&t��L4��5��+`��`NM���v���d1���~�G��W�B��2�r�Wt)K���,,
4"�h�0�A�H��Q�/xeF�3�|z�aM+X�KLVb�D�H_X]��S�Z�a��!�2��$$fs�	gtۊ	�,��,����[�T���G¿��>i�Z�>�~ ��l-����+���n�_� ��Ū����fö6KB�/Zt�s������O�����#P�W�����	�����,��we�]#,�.)&��uk��F�Ğ�K���rkM��L�`���	Th�8��I��JL���`p9�:��}�ǿ0k�ustk��bƙ�,�zY $OyG6|�Ǉ�����MF@�]��*�g����خU�S���S�4����d9��Ź��mD�n���n�U���s�APi�Ie��+k��,���J��wUK��#��*SЉ�Ȣ#�] C.ku�R�ۄ ���$� ����ԚVfם;0bJ|�<m<w��[U���U�uB��Dώ�MV�`�8��R_k^�e:��ʝ�:7�oo��D�������(�� ����1�ύ'��C�*�C�.�Λ����E����.Y�6Dc���os%?S.�)��+�&����lY\�&�@�b�f�BgeN+*��V��O5O+8���g�SL�5�HI�0�|�o��]�;��a�K�+�-������R}M��+f�f�����fk�Юr`,����j�}�R�i�(%����W�0Kh��D1y��y�YQX�O��A�LFe�~�8ƻ�c���g�o�e��zm�adR��Ɨ(Cֶ�&r�j�\]*8�_��*�8�33��á���Ae�f��v�������� ':³c��㲗W�N@�;�/�V�KN���{�m;�&k�Lݥ�����oz���V�!]��|+ӭ�s��F١�[
;�_��$���?e�xu"�3��w�'�q�C�e��>=e9Fdg$��6�EY���\��a��(L���k���1mK�މ��̠z�i��ͤ: �e�y<�S��b�,:à��Q��l�ՐO�<j���$B�gw	���0Y���[���q<$%˃���.v葟췜h��sӽ��������S\&y#��<	����D�SYE㎏���F�W���Nqm{Y�GĦB:s`��б�5��2�S�閱]
.���dR��1�
ߵʯ�?Wz�
ҔV �8JN�=�Q��<����.fł�`��g�S��<�;��n���v��兕�#A��mn�a}�K;$}�4�y[�P㎔���?l�Y�Q�	�n�#�ol �9�T���ɱ��<]Y�eM�5�[ϊ�ڲ@M-�~'���_M��n�%�!� g�l3���䷐7=|d�mQ	�w��Y,�g��0�
��+>����o�w���W!�Je��l���,�q\3�>�N�6&[�R����̦�o]Am:�O%��ÿ���LT�+�sQ3�,N$V,�&}�������f"�G����_��O�ZE@��5z�wSDW��,��}�
G�b��\T4��#��ʉ�Cό�x��Qt��o�X�ز&Ő�E;7[�K����m�� Ŵ�''���ցP�l���0S�K��Χ��I�ig�];��J��ar�*�1�d�@����`�5谀�/Y��eb�)�����P��i���e��I����U߫&8�0���CI��w-]��%C���t� 2��	��n�N���{քU���-_\+�q��<�������Z@t4aI���S�%�i�<��c]tV��G�� $0L5�0�/0��`څ���]$��r*�tT��ATYY{�C�	�<���'�:�)˵�C�`����6/�k�*��=���(�?�Kl�q��y�U�*�$�c�~ʀn��H�u�J�i��np ���
p�bRM&7~9��# ��!jl����F gB8�|�}�s�u�����pDrDPw�H��5;?���5uO�~⊁��߱���`���e�z�=��}F�cdE/��K)4
��q9=�^+����7,��Z�0O�qaY�p�j�}����H��;��h+ނ:r�Q��N ��j$	WA���{�	�a�/("1 _�P��w���g��:��S�mYbmzz��#^��Z�g�jWM�ܟ��lr������	Q�����K���)=8�P����@[Q�3�1^���P�'hS(%OՌ��+3�桟��9��P�/���հ�6�
�+P>�9��-��7��Z���W����4H/�$�y���4�Yv>���>�9@4�U/���AJQ;p��?L)��4�+H~WEэ�R'��dNLˎU���f����u�$�����rs����X|/����i�^�>���5h���/����6�⇬�{鿥8՗���܀�+��]&�I�á�<!b)\��2�'�E�\I�:$q&��K@��2UP��
�4�F��f	VҮW	?�Z<�Ie�Px5��>3�ZB񴌨 cDE��� 8��s��������%!PD�|Gj�h�#v����d5L���Zb�����$wR�=�`��P���ˬ)?ڬ��_]���xkN��f��{��U�r��ϳ���h�<��YW˅���`��b$��H6���E��y��Y�d7�#Ң��%�Mf�p��P��lt�2:�]' DH��h�%��Q�9��o�`����x���% �
��䓡W�	�Խ����Q��^�鎙�\ԚC�@3�s��[(Ԭ ��d���ӓ�	��(��Z�5�8�Xm0����KM�l3����-�R��&���v_�]هL Bd�d}K��r5&���C٣���$�̼v�������E����t���:��;�����ˈ=��.���ڧW\m�� T���a�!�Ls"m�fud��[!/M��Sm��O�8IFϤj[-�<XMԻ6O���Nm�ۊB�j��!�,0�j!t4�+�ta�%\[���Cj��7n��S�Ӈ��?>����gt�g_�>)��ԝƣ�~�f� aei������jq+8�<T~b�M�'Hw��dH��R��	2V:�f�_tAbɐ��7�̑a]Q5����C���]\wX��6��^��x��fb���%Q3�sK6��_�*�Z\��[#���Ti��\��<T�h�R~��e�,)b�)�}�F�*vUi�a��17��v���F�|`H��А�C�FĢr3�vC��C[�+�	x��]P�D��6O���V��[��m�X��M�6U�*HK�)^\�r�#����2�}��y�U�8�B��ꮒiC�Q�_�/��fĂq��U&��ډm��l��Ofʄ�
w��c&��^�mH=`��M���ݠ,�$�����k�]r%./��z����̈��Hq�v�C���'��a�6gO�y�ǜ��6TB]sy��=�%�b����LV�5��K'����=�X?���s76Dr�z�3��C@��H���b��t�/�붶5�F�C�賓�3���J��-)���.ʞNlUo��&hZ.�n���'�h���;�- r�g{�j`x�m��fV�N��8/���J�l�B�j�Y�־��ʪ0x�@���(�=kf:�-+�$�k6~ 0<�g�m=,y��(Z+q�)��+{���o߬}�X`p���uUWr�
GH�O�p�˜�K)1�	���Q!lUUP���^3p4=�,{ǆ��˺�@g��9�v�B�עm��� �w�w�k�.u��>�uZm��"������+[ 9����L�]��Y�J<5��âb5�����@�`��*Y�~�{� �d���Չ�Pz��'��Uk���}���t���a|]�˪GN[�Q(�`�Q�I���Ǯ@�Y6١����Q^�����E,�[�@�J��J������0?�*h�������s�����Y�7�N���١��?♩S���9Kc���*�8*)v���&%}�$�K��iM*�8BNe]Ia��i�F�qu���,@�Z�m֭���^R�w�"��W�i�����9b��o77Z1�;��	[�Nu�\ӡx�[
�P�&��GN��̽�o>�뎎�޵<+�Hk	7��>%��hR�O���?pt����Q��.�.n���`
��Rn
�Hm�YD��q�v�D�Pmn��y؎��S��kp�&Lq��= "��_������{3�q�:�A�&ݳ��j�B��
/Qe
ކ��Ӭ���+��ohAJ��	���$���l��zv�|�j�_�C���Ɲ?VI�(݄H��x��s>�[ǵ�$4l=�'����.;gڣI\���{�忬#�c;^�&0ʡZ��� ����JnΆ~$ۯ�"i����T�2��3�ԑ��ҿN��������O°�PJx��휵�×�t8a�H-M�細f�6�۱��g�`_,�6�3!����	j`.�HTgU23��J��Q"ckE�!5L���<��`0�s�(?gG��\��Ik5v4�R��� ���	���&!��W�/spQ���\�c^q�)��u���,/���]�<�p]t��ʻS������? �=6����K}��X�0j����oJC�r�SZ��B ��~pO�{aX��Z�g��(DW����H)Ǌ���>N�u^��o8����"�ɵ$ꍛ���er<�&�����K����U *�0�`@Х�=Dx!�G�~��w�%1X[B�L0i9�GI�y�lJ�$�*0oV�����Nvُh�c�ٳ��%	���e�5����V�Ҷ������,שpK���Z�g.w�d?5.���9�Z\�X�r�P��e#}�s�i�Y[�B�H�]51��"���+}Q�B�b�SWDµ`A1s���,}�:�c��������jjf�5JH���4!G�3�+Q��������t�Q~�GE,?�GF�U��=J���5l��)Q���v-F>,~<S`�a�� �C�s���Ql����,�Z�KV}����L�[�Nr���S���z���r�����f�Z��d��|�$��L7j���T��	S�N�I���@�;�����C����J��݀��m�d��8x �(���:0��17) ��A8Xm��|>����I�l��4F�-�cYh{B�� ɖ�j���t5�"��[~y���k
��}^R�(+���<}X�c� AP��<М�N����cd���Em#"	k,Jz���x���Ҳ�%od]$,8�˥��6����bI�e�Y(,���e��&�eqt�6���H�o�%�IX[�*߸0�9��9��;"�T��A.]v�ɟ��cPk[0����*pg�_s� �� : i����z�D��iRJ�.��-C	���>1}?�bS�UT���!Q�oR��?&�@1d�a�2�^^��
b�)3R؍{S,�=�evy�\?��
��-�c��%�*��vT6]��j7b��PN�Ǽv�M^��ZjJa�S�-a������=s�cA�zCL)�A�K�bwډ�ͥ�w���{%�a�Zy~M�NĨ�^�;�h
B�P����TCZ�w�ໝ�#�.��_��o���ݏC���E���U���#'m��r%n�ΥB�^�y��JT�vЫ�+�?��r�#u|��ݴ�ܷg�5Y.u��?�	����>�>P��;����4�y�m�	i����2����-\>8?���r��,7�`E.Y2�r\7�O��J��V�n���ba���rZ-�b�'zϸ�Gs�g8��EyfV�L����e�,s��@ؕ������c>�2�n�{�A&F�'�3>�g��Y�H*-�u��ܐ��&��\�uU�l���$�o;:�si#��3�Kbc�"[[v�ɌK�z����=\�� W��Mq	���h��1�uD���@+?\ � �������?�n��� fg�7��TW8j�xP�j�I``k��7�ǾkL�7}�� �&�\�?CE�����fG���t�E09�y5Fk.�MV�Tb��Z�=ct�O�<i"_J�Q�н���i�*��x��;Us���^����#<�a�I��;�9��}V����j������������}��<��̺�B��DVY����u
��N�7ꮺX���Th��Z'�˷�|�ʦj�KRiF�LŅ�v�1�M^��v�A��f����;���ŶK�np������?��f��K���A,b@�,�����4<
��w���XQf���@�Io�ZA��KhV֓��_
k�k%-.՚ v���I�Wh��<�b�W���('tR@����=cn��s�`�D��w�Dʒ�F���+�t+�[�JT	��`g�.Qi^&>� �xe�&N����{Z�Q5G�߮o�e��o��|���H��0���Wo���E�-/BպNS7N�˼�MT 9��2��.ų%Q{�V�|��r�ֲ޵�����,HƠ�� 0ޅoG��U���ɿ�7�������P�R>_��eGK��م���������3��Z�z~��ڦqK
4���@�'u�X�
�9��,��9�	��~s�7=��A�����+C�ـ׈4RN�]c}����k� l׺Y���VKcX@��~S5L<���@uV�T�;�g��{�h�	��Gs+�E9�'�r[}��1�`��`r��Ӎ�����Y��2^g�� 2��`�V-��Ӥ�Y�J�\Iz���/�<��q�[�����*<��QvQeg��8\����0��xs#�Oδ��mF����չj�&˻}Ld�[	̳j����LO��>�ۤ�S9�����n �~rI7��:|�Մ-�ʔND��7��t8Ŭ�YA������$1��_�qf!b�-�̩�B� ZJмs9����U��Z`��W�<����J���q�I�SD�%�$P���Q�,p�$�#lفO=jY��7���9s��.c���פo�Z-j�&������o���7��6���[���o��?݀5g��Ӭ�6�J^FS�J5��8s��M}`c�xWd�����}&lu5�܄��R��&�N������)�� AB��<��2ۥ�������L��aIZ�h�n��Έ�������s^���h��W~`��F�-%:}�m�y8�A/���Z*ޫF��w�q���,���B�փ�/?��̍mE
N���BfI'����R`eAkf��b�]��2��-���9��G��JRI����W<���Qz��+��2~�&�O�LY��?<�tt�|앣IpX잹�����1�A�7c�D���s�<�2 ��mpnR�t����?;�`�Һ/^�ct��/w�Lz��4%LŃ�� K}��cO�����1r�2Lʃ��i������,i|{������23������rP�ٯ���#\g��=P�P+�m�ie���f��Np)�
lBV7�Cޟ�Zӑ7	|l�*c���q�Pk1�����9��k��)K�D��p>0;�������<Ah!U`��0�����oQ��h}��fˢ�=����U�}��b�.�z�o�A��y����N�Q���D�L+�J�+�v��h1�-[n�Y�s�/'N�k(<�����4�CS3U�LﰌJx�ڐ�_�O�X�ф���1P�eL���� �<�Lqu
�T�8=A4!��% g��cd^�qv�h�W���i���\�-iJѡ����e|a��qX�Zzȧ�0��n�Z��IWVDIV�CV0�j�<�#������� �`;d�cwg����I~ά1�5G7SCļqv�y��#//�+���74vx�]�ާ�H��������$�9��]T��-�u�d�����~���S{�`�(�د���:��y��{D)	�K��*�2��4��*۬K�yL�ow8*?���SE�O���(�~c~B�v�nէa;�O*!C�qn@7)^�\K�����Nh��ɧ����;��&SǞ)�@{�K��נ�!�4^���v����-M�L�3�pqHd�����zf�覜;i����ZU�vP��{�y��	*�u��������w�{�E��>4�x��4�n[M�:Ơ����;̼�+�ПL��G%h���F=��/�®vQ�e��hp55ɭ@�/YuO������㞱jK7A�	����xb_F��o����j���k�t�~F��P)�t{:]��`+�p>��@�]h��3����W�k*�3m�y=��F�u�M��r��_�(�1ȃN؟;��N�l(�fK�*"�*����X��#R��
���q\����yGC!L��hI��8���QӕK�A�W�,�cA*5��wgsH{5�jt��	#�5�%�0\�<$p�P�)z9�Ɠ��aIA�M}��#���ֺ��7|"u�a�E��t�Vҩ����+6?|�R�pR� ���"%/w�8Lc�n���E����Z�g�b�cD�snk&I�G@dIUt�Ɛ�����a\XC���dࢼ��U�0YS��9�
�.�Ӭ�d�s0��뀌��Mn�>�9ac2���0�7R��V��(�I����d�`�v4���h)q��#��V��˾K��z����DĐ]����Q��=0����&F���C��o.e�)=[�b.`'�.O��^%I�6��T���:�b�%5\�P�=�0�%��_��7�u�WC��y[FX��� �?SuO!F��]����P�*���oD���[W٢[#�7�����~�x��l�);�L���[h[�+�	;.�Z]���c�0�e��ݽ,a�rk[�2����WK�� �Υ�c�k|2��Ωm`p=d
⬀�5�_c�/�ތ�h0�Pu�7x7nexz��o��v	�l�0-�i�K�ݸ�D�
�V�>��3um��nqB#+H�u&\�d?hV������N��J��[��wo���x�3O�	�nx�/��A� �`��d���6Dܔ�k),�2�9� F��L��FSu���Y�h�q�e`'�ab��˂�+v��s���0�xJN��?4�?6Q�'<>yp�%�9����ь��t�Ey(�H�)482� �>Θv��3�_ k��}�C�Ɵ	\D�إ1��0���TN�jyB/�Z4tP"�(w�O�v��Hwo��?��M���<�`d$��j\x�g�+#��L�G�`z�M�2�/�2���^�F��@ӕ������Q���pq�Ú�ؓs?Q� ]Oz���O\�(�p2�"��%8�R�a?�)̈g�1;7bW#���%bl�<T9���t���)��E ���m�Y���N��%[ 3Y���\����ˣy�B��"J#J��'�=(L��0~ʨ�/XB���n�p���/�s��z�%Iѳ�����M+>W"���Di݌��c�.;޵��h���+7���U��	��x�D��M�8���4U+�w�!Z0p��;�>/n�OB�M���U����Vf��*o�L�&_��7�~s��������Dȝ��J;���W�60^��3�a�y�^�ii�.��I�Q�]ԘT.����`�� �X"$��6*�L� �>,�"�#� �R�4*�J�çE���(�]h��'��"��]����e��x�(�Еt`r��S���F��a����X����xJ֪q��7�B������N�Ϗ�ݘ��F�B̗����z \f�[��`6n��9��a�u���4�%�_P���V��g����Wg�(��a`S\c���������P��b��6J)ltL��RL�F�1�@8>x1Տ1?YV� ���@��Q��R��+�ىJ�F�"�)���!�Y�3���+s;���!��_�y� �1 JtJ��n�'pT�&��f���c��DY�\��"���׊�ߎX7��W;M~+P̞�'~&f��̿ud, Gk���b��٥�k��F�{�����*���3�������L�DSo{��Gk��C/"e����Ɛ��^}%k�T">�y$9����#gD�V�͡�o�?��Ȩ	�x�bSg���MD���NF�n����U��D�*'/��?H�,{+yd�Tbޤ��S+�Kŭ�1
&c6��]7h��	��ʍ8QMU��ӯ�#���f��o��[Y4�w�-�i�Mf��uGm:�<���h�?�e�I}�!@���L�THM�U֑ž���z���I�T`�W*�?C��k�jH�v
�^������%JѦ(�8�D�tn�/k��tѩ�g :Ն��y�O=�����ĸ���I5��h�k�B-򥘆\w;<?���٣g" ՜�����S��0�wSb%Ӷ>ԑ1S�CM�~��	����8�Z'�K���~����TT�ǩ�������=6��TB����qU��R=���P�+��\�>Y$�;i3]����T�����i��̝��߻޾a������mf��5�+J�	ET�5���MGN�$��Jr��Qq=@N�M��)�/MK4��� ����LS�"kR�5�4��W[���#<\��E���$�ѣ��lX���$/��%ĉ���"Υ�X���]"��Ș�MR[I�s�P����K�}��>�]����|5]P��4T�d�N�h�l9U:}���Bd�ctmZ���h��UnA;��O�(��UZ�Ǿ����㴒�ݑ7�ǍP��d���x�-q�e��Lk*�����g:a�N�"����]\�
]lE�L��h��P��x�Ma����Aqd�~Y�����f���"싼9B���I��#5͒���E�,o�m�ۈ'%���L���]Bx�� �"�����/��lܝ�5�� �XP>�����_d��GR��\�{���_�� бg�;z��V���*䆞U�k�s�z�Fծ�5�fk�W��2��X㛂��!�>uM�>��ꡄ��eMU�A���sh���*�!?R{0�urO���ƾ��Mp���'e�!
_>�+i,� �~U'h�5N�d�����S��I8�����MLz߼ S:I��Q��g:�pH�T8�*�|��Q���̂��"�[�!B1�4Q�1,:M� sH}�u�I�D�8�M-�X�4��~Z�+yQ��Yj�u.T:�C0���lDd�z��mR�2	�y]�l��Xv҉�/�7sgs�y� �V:��n��tS��X���]��D]�\�H�-��=͡��T,�|k!9��)Ĥ*��¨���](a��A�����\ɠu��lw:0�*�ۋ	��ǯA�şt�(���WF� �Q��_Y��Hv^!�"��������R�.@�E �\��`�1����ܵ��|b�
�cx�g��� ��cPܭU1=�X��NO��c*��>��ٟϚ��e�p4��&�� qO��i��" �~��
~��$���h�f�� 5�;	RQ�|�cX�o|d�f63���q8˴���1�=�	j%�#k:/�����$|�囨V�Z������J�f}�J�uר[�D��v����4���	xD	�b�7A^l�H5�c� ���N������p�+�I2
�؛�E03!���>96U�(U��:��OԔ� -v�*_��:�V��/��>��qi�N5|ׅΟ�zF�2= y��h�e�VbPu�\�j���s��b�Ai���dG][ߌ���h# ���B{r�)� �����\]��A��8�@��^_��
�"z�0F�-@#׏G�v�!��s_��OѠ����o��K�Q��r<�6�[�uZ-s�S(�],�[%f@�������؆�w�a ��`��6�U^+�2>�D�,�dEKZ���}ml����x��M����r��	)�&�3j�f�\��lbГЦ�1�|Y�~#o���Ąc���E!����)��k�)���&Ɣң�#rU��E�4���`�<_��B�HRV�x9N��LCӉI+�'��Y��س��Gvg�{����5�'PtH^e$������.�i����d��5���t�$&���Y�8"Ֆ��(�$�: � FU�oF����U�(�n&oc�>J�1���y9N��?�L��O�W�
w ]?�P��Y���͠W~�.�(D 9���e?��IcD�۪!~��?�ޖ�s#�SD'�`�vvD݂��q	�w�O�F��p��wv$�sK�h܁dE˱}m:O��#�C84z,ej�A!���tA���I�2Ѣ���{9�^bd�52�|��)�#��6�����wi�C5]�* ���n��VJ���Q�{�Q{b
�ѯ�7��Lղ؍�Z�cY۵����}�mW�^���?���L�*ot�?����Nfɰ;�����I�iȔ���y\ps�=e<�C����zz�ٮ��K��3�D�y�D�+<�e�������q�Ľ"ء����W�'|"�؁�	}V���OB��m�|�]H��ru�-ƨ� $~�&�(|>>&J�D	��V��{+��V��΂�#�X/դx��}��c�m��x����ȃ����1�Wvw����xǂ�&�"����p+����/���q���$�g#X�+�2�)
�q^��T�k����S�������P,ҥ�v`�d���a�@I����W�n�7����(��k
��G�V�q/ju�e�j���1�������s�y�yhi1����t��fo��;��R�����4e稊ϲn�=$�`���~�Ep�B '�xג?"�z]� �}�ӌ-��j��&vL��J��Z�.�\I����I	�N2H��KtN��U��ր��vEf��6��٤����cRJ�`'Ԇ���N]��ŷ+ZVM���@���C����}mG2B���s�z��~kԨ��;�e�[��`{�,�aAs�c���%���mrb������T���2��%�;I%�����E7Y◃�{z���nj覃  G���	��v���v��;H����
�i�zxBpŖž�N�U<�q�1Y6�.�&�&��h�0`�"MΗ9w�Iݯ	r�y���d��z���  ��a3��=�����Y�nv��*aP)F�4�W�Vg>ֲ�	��	E@I���^��*����4�]dԕ�L��$Oy�Xd���]�̂�� w��J�b��������D���mfȣX��n*��}�x�!�[���{m٫�B%�, ���;B�[H�]C[zd�\�
mS��4�F��* \A	C��ѵ��z���WJQ��i���
��,���m�ǽ����%�18HQ�ŵ�����A1ꖦU��8�,ң��{��gj������������|�����Jl�R1�2�7��	�~�f�M��.A����Z7G�bsZ�_���HL��Rl� K�v$G��d�֡~V0~v l�T�^o��ј���Ds=�B���"���h��-�����- 7#�pڭq�E��7�l��>4���/��N\TYY+�����T��u�j�5(�;C�*�6S?�RX���q
�.t�V���t��)Eˡ��P5\�j���?�j��*7] �&�Q0���f`�og8
�	� �o��՚�~��iٵ�mx���7XS�~3�ǻ�tS�-�Y���;����7����չݢs�k���ՙ��e��Nw*+��Xp��2T�v��Z*�;�����ap�5�\���9\u�S�W����~(#��ج�y�,�g��>���g�m��u���>C���|B�N�����,4������DrDL0ڠ���ś��ʎ�O^8�?]���3ȵ�@"�,K�����������"I�p�ne3|C���]��F�vY���H��H)��-�9fu�\��NLŽN�ܧ�����<���{�q�
�2R�i���au2��Ґ=��de���T@3|��v��&��2�:�t��\��g0GX^q���8J�KG�-|[7�Ƙ���B���!�0Ԁ�mG�3�3\$g2�[ws�k�$ =�w7��xe';�MST��OFs�<�BX�9\��ܾ=ni�����.���9P:)�1��O���9+n
p�E�/N������}ش�&�3;G�:s�!H��ͬ�|\'Z��y�rf�8���/��NK,3��8�H��e�5�����+���	�<����ז���(�R|t�hZ��ä���Z1�n�c�0-\��z���?p�ʧ:�����َ���wF�%��K�/܏����n�~������5^��I�F��:�=6�2t�TV� �ω��O�!�I�'�MhѨ�JK�J5��(�iaxB�z&5�U���Tm�ϟmk���G(M�D ��~�͠�uN���?�o��=aW��/Opٱp�� ��Is��0�br���]7��
FpÍ'�I��+���ͺ�F�%+�$Z�[	@�����j��ynm�RY]����l��u~���~d�J��?5�-�y���p��T͉GY�䖜�q��ٙ���P��zN�˵�� 0�4���򏢚��\�]�ѸܩZp�R8u��0�[ˀ�i�^�)D3X�BX�����|jpAg�x�/�{�Vx�g�k+}��Oa��ج `�N:WC�U��Nߊ0�-P��-��Qo���r�Ze>��i�>Lsr�ϴ��KT%�L�"ӠK��D��R�=��sn?KF>shS:��r��C#�I��o������Uw�l�o��tx�y��}m�.��O�
�LcاB�Q-�޽�6���|E-�D3�iRIs����眥l��}G{+R�E�ׅ�P������Q-}��9B^^A��q�� �H~�^?�J���K���Պ]���Ѷ�����?�����'��m���u��z����A��ᔥ17=<�1�8�v݀���S�wH{0w�3�8"�՘_�ˑ��7"�s�s0�'O��OM��%�פù~����7-G@�׉+!��;���nj��B�?�t����9��h�"���_}��AfD�-q�wpf��˂^9������s�Xj�p�WS�$(�e2索�p�jՐ���L��֙��X���9��K"��A!ݍ΂�9�5���l
�����u~	o�VPE�k��R<%`��O��s��a�t}�A�r��Ts�XO����܍bgQ�H���B���T��o+�7�BN�K`��O��XU���ϕ�Pїly�8Tx)J!��2ԥ��/�j��&[ύ�w#�h+/�hs�W]��\�	�t�7a ɡ�nh��$Јxg.B��z�jr��ϮW��w҉x���	���\�?�W��l-��67����~�R��6z)M���O}���C��~�t@����!�Մ#`סS}��š1B�:�m+�*�M���og��F?�����j#���l^�9�Ȣ"<A�{F��?r�ح��xv�]��}Ռ�7#�������#b��Wt}�j6�@�ܧ8��fwͤ���H˺� ��֚wd��6.��Kd�g��.1�2��z�u�֙��3�y#r�kꈾN�̈́�8j	eh�\����t&ن��)H

Q���e|)=;��0������7��<#�GZ_!�i���#��	h�+x^�;�?�A�1I�Uxpv��s�������tS���^����q�1'v(4�~�"q�F���T�	��+��jnVS��G��ud.o�Y�r�ŀ�7���D�����Y�p!K�"临�Ȏw��\�AnE6F),f\U��Tݟ<Y���^w�ӌ��b�t�P��?Px]��s�Xp��Q+�-U}��Q#�r$딣UC�	zF٘ j4�#�� ��OL��E.��c�y)#�rZ�	�'�*�^�:Pi(m�=��T��a�������BNBC�)�9ޏ��J2�T�ߕh��9�J
��7���S��u4��_6=r�� ���5-�_�R�d:�4j�9�� W#��Ȗ�.�T^��A���Hb�5���$,Eʵ���lZ\_2�!)�������P���<����^"O]�TN�ӷ��ooEA�9��r��Z�`�Q�\儤��`\�E
7F������`���k�3f��.���Xx#�f�k9�sH�&B@dLkqF b1{�Óc��hɯ(s9q�3g�}��4���܆��繅"�@���s�ݭoX�����<�� Y=ꨔ��t6iѽQ����1Fb��T�_�س��I%�cx�@8sE�q�� �1���S��{=m�Z������B��4��XMĮ]v����1�_��(z|��7^�ԣٗ� ��	+X{%��u��&t���@h�O����S�M(�CJ�2&��4���W�s�����/���8�1�ٕIPh̥�1�u���� �����tF`�7!ʍ���D_���Gu�yK��Б��NP`݀�)gLo���F�a�M�uC�,�m����ݑ03�G�D��ۊٶ5e /uD-E��h��J������Mw>i\��h��<=iIW`����<�cl��$~�Ϯ�F;�yQ�*^�C�<|���R�';R�lf��gů�4.�u�4�8�A��qhԱ�|}�2ע���X��Xl$��/�@<��r�����|36.Sa[g�e����hS�A���|r;��O�$�8ꌦx���"���Q�`+)s���c`����'��Y�U\>=�f�3����^A�a{��G+�A� ��,!�M1�j`���K��cO��EX̡@M���g���.�����%��x�oPe�;N� צU�9 @6뉥h'�͐\�ܚ8Xf�9�r��:�;��?��n���)
T*���v���Hr4۵�C����̐/��, ���|��DߴM�қ���*�4�r�4�b�^)q�+ni�D�B:�N��^Ċ͎�ԈaM�>�~���a��HM�;��*Ȟ��+�Q�WQk����[�AͶ���@u[�RF��:��eu|�>Z����1�K����3%bg���;Ջ� "�<k��`��tK��~cж�¹��>%�=>.�m��{W^�N�:��ZH�
�,6۱6k���c>J���̥o�QC��7�����	E�q���*A�?.���6G����D4x�U?E��������� F܀���La��7U�ӘN�9���3@�P��ѭ�J�߶�'�;�����Q�5j��،E=�y�C�V�]dU���d�һ%K���d��]����@I���q��c=�	fۗ�)h�zAϩI�õG��X[a��J��zb:=Y���������g |Ղ=%��5X@����9M�xK�\�/AI�b��Ԡ�
(- ?G�:G�N<�_
��wS?9,T�b~�0�;�5�����Z���a�To(�f=�hulSR���B(I�N.�y��kY�\E���S��51oNp�cW�㣈XڢK4�/��c5�.+`կ�����)8X��\'F�m��5��l^a�Q�F�P�C�K�?����j_1���pE9+��c
��[������!p��7�ip����wߋ��D��V q5?eC67 ����_S8��O
��'n��۱N�|�k�!�ÛV�B2�iz�'��D�]�t�Z��]vNa�,�/���A61m�WX���)jՙI͟���#������$*�g�V-�T�n�����%�	I�3���@�e��)$q�p��/����PfO�z=wJO������v�4�N�(�p# ��B�ܨ��k'�EǵN����_ݽ�a�",ť�s����)蓮�i�!��+7�(k_��նF�K�g�g�(XKZp��;��TB(�u&�,��B��C<AA�B� z����J��ㄍ�`�N]���#tMY�@6�+76�O�T��|�#�����`�K>�tz@M��GO�|!���_ċg.vY]n�J�(�QXR����[`�aT��{�������}l��9��1|�X�WK�84��9�s7�jć�x+�-��ɲ�2���~~�i�dd	���U�g%����*p���t��$�c���?^��	��P�!�#���J��I�TƔ��h��w�t��n�f���
�3B�V���	�~t�|��PMڽx���ԕk9�X�

[)R=$v}�V����$G�Nն��V�������E���7��h4*�K��=2�*މ�j�D�SYy��+fڏ:<��f�E��/�L}��������:�#�D�7�ck������*��HV`�)��4�#��:|�?��_�}��m�@!϶8�XfC��ȼf����q�" ��c����q��ގ4����]=��KQ��S*�s�ı���N2@����ަ�֧%�gb,�J�۬�f7qB�
s��j�nm^9}�3ĳ��E�B. ٶ�����m��,|A��ʇ���}#[�M���s����}�j����x��'+�C�C^2�C u��S�v1�{ғe�-��ЅJ�Z>S�����[M*����ѿ�&Q�qM��ǡA!N�����s"rOMJ��� ����K�V[��!CN�]C�:��WE:tf��,�1:D��e���3�%΄k~�K�o�P���i���F����lk��_?���N�B�Ȏ���Ҵ%�Ys��t��DV�£F��3[���ױ�E��b��N \ӖPH���yއea��]l�Y��*��x�:.g�$�Ң��sh��Ll���!��,��_����=t�/��f]ƍ��S��@܃��%7:���:�N�6�a�f@9:2�������[I"1�z"
5��$0"<�/�v-`A�"����ȑI�Qr~8n���ˏԛf�xI(\�������tcP=�H���Vwʜ/����
1o�Z?\d	~TL@bK|[C�:��$L�0{�i�]�%u6�����5+`X����T�w({m�����=�ϥ��	J�&�5���32kg�Uѻ�}�<���+�'��Qk�܄`�4R�0}U�/E%�m�š�{����&*���9�Dɨ�D�j"��
\[�D?���rX�ò#I��Q@����߷��qe	��:RV����W�����X�n`����#j��ѳ�Ճ�fR���B���B���X ]�����ux�(��Ng����M�ZL�]k��a��r=;��
8~�,gV��Ƚ<@�0��ĆQLm^�<^�jq4@&����(2�b����m��<�a�_gܿ�"�&tH��6�SL�4�	Q�Z�G�b��(�i4�O�ET�F��ܩtB��ER|cޛ,���f��m|��6����ʮ�	����*,�w՚fGyif>��Vn)	��q����7��9����4�����4�v��TI�����U���N��	�t*e D�K�`�Ud�;YN8{�%��f������۟*d���֮���_DX5��HO��/Q��ϟ�1�(�3�>׋����I��I�&g�b�O��ѫ~Բ
����boO1I@�1pF^��}��P����Lu��.�'���I��Sۉ32���yG�0��xa��0��yB�P���3���b%�Z�K���M��R� '_���2��5E�����79]��B��Ċ֐'�,_����QV�4K$	'�h���R�U}�T5�]��kd�����~.Ι?��}=�#�����Д�?�~�v�M'`I��\��F��2vL�|x����#6�}v�d�E?��C"!Fi1�!�Z��qV�nU�;gw6�l|�YT�e<Z:�[wH|��9Oi8�'���Ӝ|v��*59��,�rb��Uv/~�(����dv V�׹���\�Խ{�@G��U�\/���B�A"�#ZY�^}�A�w�o���n�g	'5�벴�=���м�/Qq��S�A�w��.N��w�0zV�ҤP�9�ew�����ۃ��:]��nfS��ț��x3����Y�}�tA���=�)w��6(�koR�@���n�� �a�)�]�uq�����&�� 
˹G)vV����.k���;��m��GRYt_�o8�� �N(�i������I1���'&
8���XA,����ً�c�Cp]���(��h�oX��tr�'�Ӈ���(�m���	����u��!�$S����͖�L~�|Ɗ�d���1z����~G[b#��ُ=t(0�d�]*J�\0|�~2�1�o�,iЯ�a6$4�M+H�l�D�H5����e�D���5.+�g~%ƚ��JwB�`�[%�]v�z��'!@aUX7�*����1!����&Uѯ��|`3����I���y�*i���a�$>z&ֆDi�t�-Ơ������CBx�eFu<���I��>���q��X�W�}��*�yð�� ��6�w� 9�9�'#��p�& �}rv��z$��i��`4�nB�	�֓`I����y�;3=IK;�LС�12}]��ce�x����t��@��[>2���A����Ob����d�W���X	���s��
'��о����է6��AT��LH�2Ix9�C.�r z}��Ye\L `a��l��#�Ǧ���1�gep�;����V`�A%q:M����s��}����8��}kn��ك��B{ �MǾ7���c� ���a:ky1L��,��|�r8<W��g=��Tu�K��QZ3_Ȓ�K��`�XS8pm�ߟ�d���W mF��+z��c�mE�A�$��5�Sn7���Tm���2�2������������� �Y�����~�A�����*�A��r0����H���}ہQ���m[Ÿ����	eһv�fD�Q̋�ua�W����ޮ\�D�|�gY�
��tAխ�iNl�X�H

$��lވs��e�{���G��Cq.���9`&fjd^�a�+�"@1t��9��>��,lA�cT�+$��)��H�9a՞I;��F#�57�	��+���,<�����R�<G�c=by� dG�y ��l9Jv�C��'�k�!Ib��@�4氛_e����"J�]��� ��W��}�c�3�-���0D}�t��֡���w'o0%����s��ގJ�U��v[_� ��c��O�F���K��r\�>*�\N�Z#���x��Y�6���B(���~�u!���4�������L��C� \�D��? Lݑ�ҹ�5�M##�)h���#��#{'��t���s�JG���K��Z��g�<Eb��vM�-e���g�J��L A�c�*�,4�7���xV�i"03O��}Q�V��Fa��<�m�-A��D�8�
����Ɗx�h��>�H�����"
�ć�����.20������g�ڗ|�X�)�}k4��N�u�g�[\�|Ƨ=�~��W�9�L�|�zy�u�zK��ݭ�ɽX�m�T8G�Ę��)/���#6���������\�.V4�{L�G[�DO����/��&O����y��N[������B��:��{��Q�L�+�Ng$3q��&1��N-�j	m}�7�s"��8��ʊ������}m 4*7������[���;�QχjBΣh�2�����i�C�X�CFy{'ar6�I��H���i57��Ԣh��3�+$���t�92yf��^m�ӌ��1������|�b>��Iy��D*'�疟k��~FI���p@]J��45? �Ԫg���mCG�d�2�ϓ�r/�M|�^`�z��s�4�%��lOC�K��e�&7�g6�@;��`[L�rk��3��$�$vV��jK3vs�����*Q�E����uE�c���要������QӲ�SR�r��rLWb�*�P��k@R��C�Ӓ�4�"����Ɇ��
�7p����ፃ�͇a6�D����q"p<Шj\�-���1k�t���UU1��<�BAG��Jv���?�+C�!@>�ϳ��*M4gP�:{-@3�>e�AG����B{���+*BQr�֤F��=}�!)%�b�H�V�,O~ w���䁙�f6��z���O/Y�G���+q�_.NjG���mүW�^խ�oݵ啈{�^�� ����/* ~�>��5�fs2;�*�S�iT.�d~��cȞV��,s�OߖǀP�����T+?1Ew���/~�+;�P%
�Jn�9C��&112J3*L��Y`x�Ƀ�(��a
pՎ;U���J�jmֵ��Z���A� s/�η�h������HO�Ȯ�ˎ��c�s>����D�V���{��D�)|x7����YQA�ʁ���;K����/���b&�t����ߙ#�eb�y�����es4EV{�h���t���q���	�}ݼ>����U���D�[�^���a?����.Q��u��T2F� �X0Š������Ț�B�/�򃄍)�Z�9��T���1�������A��y��O�����<��Ь����l=��Lk7���_`���� ׿tw ��!#+u��o�<��=�RA��9'����iwc��vq�↎���Ee4��:s&=�o{�F�Ω4n�dk-^<��o<�hz�$�Z�j��+�0�-�%��h����W��>"?�C�۵�O%��� ����G�~Dg�Ja��^�Wۮ��ǐ�F����ғX@$ySڣ�F3��=�L�����<9��n��*8�e�{u�J�
I���K�e#b�g[l��s_��X�]Y8��o[j�
/�D!]5��Ң�L��F�M8/Į鴐��`4'\�N�A��x��^ Z�+�"`�����Q��0Yz��!ʄ��F�-vN���kF0%{���%xjDhMj���C�Ik�������Mԙ������&�$"3��m�L��q�@`L�o{�l
q�D8��%�%����_����y;A�z�ٛ��}�̈́\�+tsR&�/��W.E�1�4���Ƈ{�^"��X\Xc�֑�\!����Ys��a2V���O����x�a{�j�||����������htͿ�2�~���"W�5��� ?-&���,P�#���z�J����;i bv�����+��l��1��9�T:%}�16^m��Ԟq]y��zPY��5Z�n��֋�A_���yb�j��@1�U��gaʩFP���S{t��v���7.�T�J��4`Y����ć��@��I6�u0%���
ѳz�`Y���(Bo���^�DGǱ�� %�X( ��eЂ�dz��,&Q��?�����j�O��o;a�a`T��*��v@��=6{R�*��8)�.��J�����nx�u#�ĐX�l�`:mGF���ݣ��0
H`�b\<%'3��2S``miH�g�Y��"o��I�,��;-��Ӌ�����l���)�a�SYQ6�)�z�����2e�=~��_�]� �a��ڷ�돔�TN���C�k^3{)�Q�.��,��ou���O�_����󮷅����R���`4�^��3t���]����N�f�P�ҿ�����acਊc��`����*rm�@UG�B^X��}�Fex��6tl�oć���Ev�q�}'��U��v�D3c5<��X�y{)��Y��.����;ĸm6��'j�[���v��kj���/�v��U���(� �*��{y��8��	�u7�ճJ]�ٰM�����6�` ���g�8��ڮ��J�����_V�l�J)_NƧ�	q'ĎBP�3~����>F����xfW���/]�:[@p|J�b�~���1��Zt�C4�J�����fw���x�Q6p�53p��a\/XE\���Kn��6'>����9ZD�݈ݡ�~o^�^�����d�/���������	P��Řf��a�uq�v�u���æ�³�'���:Nz�-d',�lg���	�߄�;)��Tpn����C��g��� n�������S�.*i��|�x<3V~-�5��"��u'�"��c��)�U	<j��"�Rz����_���A��.����
՛�Q\)�o:ȃ�$��`��<��L+� nG��+��X����)�!����cR�oeB�-F6��S}m���V�h=�{��]�#g���X����.%C���4��Z��t��\ gؙ������4jgP��R��̲m���=�3��c`g�1:ş#�������	yg��f�ϯ@�Öx�W��jg_J�O��j�����l 0%����|L��8���Dg8���b_���Ln2.H橃{��#��������e�5��X˰f4�W��	�7�	��m���<�׮.�����fvCץ7X���H�������l�[b_%̮�0���t=�lf��$�{���]n�&M�7�Ԧ��,]xUK�:[Ց�f~(��Y���.z6/�y����3�]�F�SJr�z���A�;1��'�{�~�cV�FVh�2f2��*�8#N�/-���������~c՟۝Q��v�������?U�L	�%�ڝ{���o�D�����f�n�3��x�_�69��'���)T�v^���8G� �z,��5|���R�i}�(]�o��[��Q/`4Ue#i�nXS����/�c����5������3�ȡ�\٘��h�K�@K��T�C�����-H`�;��E{�%��LK���Ⱦ����C��΅�ʇ�p�Zj�'T�0ktaI7Yc�?�<��:D&�����z6���I�� ~#��M����(L�Ԗcu�d��YK �����pnz��ίG����s����$?�ގ� ���`�ID<�M���� ��$L�A��-
-���3�L8GJ���i����qg.fߦl��[J΄M���/��\��=ľD�Oy�F��|ߌf]iWR!��̆&����cm2��j�/�L7��i���՟cTZ��um=��]]���ʿ�(����
Nl��<naA���r�߈��䁡�J>�e�+0�'�5]7���H�q*���l+4Frw�|Ra^�ım_�����������+ þ��c���!X�����P�Y�)���S�Z�-5���FG���b��3�Du�(C���綠CB�F@�C4{��-�/�<Y��X�?�3 y���$@�&�(��l�y�����ۑC�7W�
�B��������£�P���8�^�=Ι���0b�����Z�a�q�Q�8�A����۾A!�wi��gխ�e�3��9��7��d�s�*̍d��e�w�Z�� 90������r,P&�K�r�V�WY�0���C(֏ps,�(x�``� ~t��U����wu�݁�G#�̛��w᫔�]�\�pV(��\2����;"�Xk��ۉf�/�A2h�������j_4�ʹY���}&��͟ґx�	��(�R�R7�1�.��G�F��_�μ�U�Q���C�ڍ��1���6�.����j�9y�-k�������l��*��o��uT�`53I���E��j�c�^-(�ͿAB��1�ؘS;ϥ��_'�O�e7��h���*�֣���0�zH|-�ˁA�$���j3iX{����d7@��i_RsG�!
Sk^E��e��P��UӶ��
���?[�.�����|>�El�F�������o �)����@{�q��� �>S
�F=v�ɤfg�����@.�k��|�jeB��>+�8d�对/�s��JLΝ�w_�P^�BF�LY�Q�6�G�ܪ�]̄ߜ9a��6W#�<�d��Zq��$�@	%�����*v�f+�@�@��4�PLG�rh�'a���r��ciMK���hۓa��#@i��m��=����?��w�[��Qc#,.Eͩ�׏��1��[Q��ِ����#����5D���H%h�ٸ��D�n�� q�����\>�#�ϕ���~�B���V�`�iOB�2P��O�ȉ� =��Q�t��РO$a����i1�����h�L_�c���?���<�􁇳r����$w
PǢ�N�2\��|%��vPΕ����Ćd,��89cp���*��:��М������Q���/�����T�/D�
�U��uC���t���b)��FK��8dOGk����󝯳�B���ݼC!����}B_�bKI��Gb���@���&�i���y��Ll6 �NPk��ŋZI�5��A�����Z�g=��{���h�t�p�Öz2�h��\�2^0$��/���m���3�bv"r%�F(�#!��+r�#~�t^����n,���QŭOIɡ(�Pp\�S��EP�q�/;5L�8���H���1�+���(��%�f�AaZ�2$��0o��4��6���~z�˺ �m2a)!Vt�����ԇ*����)�"'/�
�m��+�d'G����![Ѿ�	��:z�؛�[��[qf����'W�\w��ӈ��K|]��:h����	��ֳ�B~��8(�����8A.q��3)�|���w$8���{�~�*��ܑ��ӊ͋o�NMC��H^`�$�p������
���>�fHNLWgٔ$Ҁ�!�)6�F_t�iM��g7K<�׾��k�&{'�s��& g�8�ֱ.�Ev�{��ckw0+���Gy�p��D��6X�ţ%��Y,}��M	�Q�:&l���C@p,�e��[hX��61O�v�����.l�,����
�!\�����\�g¥�7�͗s-
��B�؎&3=�zLa
�����KT�;Rй�׎����q��P��;d(�V����0�qu��3�䁊f�gUHe�YZ�Y��[2��w��nJ�_�z'���ځ�-�~W���n� ���^��4�v/�4���Tf��b�X�����O�����u�B�Ug}��7H�ᾩM٪��6;��8�""b> ��t_���ni�c�=z('��9�5m��	��7v��	��	C)�]Q)SH����Ɠ�DK�����[[ab����~v~�U����#X�R��qv.w?�E�Qn,��r�̐�8�pL�\��%/1ϚU\K�}+��BP�2Gu��*��8zy��0�׫�����ܤ�:KW9�36��|�r�?�d����ډLd�yS��C�C���0�`�A��w�I�"������!���|�3��B)><�z��ϑc+�v/�����}[M�<ے
�����g�Vd΍���+L��6�Aj׈�����&�����RW%3d��賘%T��g�r�1�B��Y���J�E�Ţ};m�a��i�)4��.>���"��|�X���t�fâ\�g=��L;�/�:uiB8�4=- v��X�ә|S��UC�;b�rwsP�b%+�2WႪlS\a����X���p��RL*�iQt�G"�B5z�l->;��轌/�OZ�=JQP�nb�tAv�Y�0�y~����J�G{h]�}�[��B�N�>��}�����-�ӆ� �����q=<煉�ܠX�Ws��k1�� ?&�B�4��{ۆܼ�ҌX5�(/6���:Gf��(ձ���X1*��bᱡ�9�����.q2�\<�:����bm"���!]��6	�LUqxM1�$.��􃒒��]3���AK�2�3=�4�@٦��$s����66��*WѱoA�XJ�u1/�EyK��i�Emg�M�
K�WHM]��+R����/g��� ���]�75/�K��ȧ�B��ۜ@5]r��%�*�[��5��5ƒC[^+�+o2�{4��b�A�� ���v��9!D��w?�1����q-0��+�L͟=YY�Y����u":ˆG���k1��׮?�on��hK���E�qEު@K
�87�-�a������3yc_,M��������_�F�˦��c�5�K��߹c�s���y*�"sͣ�����h�;�ޮ�e�Jx��N�5������7i��-��P�R�G��ԚϜ�A�����eq+b�鷤���@\���s_s�M�.<��~}���C}��H�ĉ𱙕S�͐���W6JD��~��C�l"+Y5�$ΔV���Y�yrtP;elޔ-���b 2X�u|.����|��X�Ug��� ��#p��=i6���$/k�X��a*�zs�ڤ���e�s�m���h���Y��#s�z+�c�{�ѣ$�vem��oM/��\�e�#������_��9e��23��I�~H�۪.\俶PxC����[��~��/k��ڝR+\��`E��M�͌]A�)�:!r3�����a�������9qq�z������m�kX��Vk}WOj&U�B�dپRyU��&y��zT@���lZ�~�V�ē��W����m%�B��q`�Bo���_O�{��qj� Lq]�{�B���~3x������F�ԋ^Y�4J�_X}�9f���az��}�w�L��pŌy�_QFG��벇��֨Ñ�9�g���fE���H��K��!\��m��=�Y�kI��L �荡�۳�&�ث��ǰ������s����덻����	���1�U�Ȕ���˽QXJ
}Ox\���W/�HO��)wbA�l�nF�
`x�lg*x��~��6�I�I�"F]�n�X�
{a�V&6BmU�鲁&E�i��<���*V��^]aB��1�c�KM�a���m��P��#3�gkW9$t?ʖ1�
�@�C�)~x���Oq���ۧ0%q� ڝ��-گ�YRXD4�,`��T��^�4��GY"(U!Y��5��#§]��d8�L�Y�ZA�e�jYp���H�yM�Y�z�i��嬉/t�]��
N}ˎ���6�g�1�f\=1�k\O�҂�o
\��,Iw�u&ȅ=Yz�Y"�y�o3�֛��=�Q�����}0�?_r�!l �뾨�^<�Rs�x?:��=�ꛞH�]Y=7]Ȍ�R5Od^g�W�+�A���jz�O�í��Y��o
��t�G�*�����A�^=�y
���Xə����۩�0CV���%]�J��Q� �F��w��\�aQ��PW�J�ԫ�p�lr�Ý}�1�n�t�>�-�.�h�����/��&Wm������ ���nwL��UۨCY0�w�p�)��J�h\�8�B�=�:��ٜ<5e�C�T2r�^����.�]�l�X+�d��v��&�ɢ`�^��M*fI�q|<y�Hg�֯���E�����M�0��V��	���4S:�q����:<	h��9o�	M��?tKD�e=��m�UI�d#�QL��m5+3&��"9�0|�VU�6M�-ݯ��"��Z�Vs��}W�F�ռ6+:�Q��μq,���]ů��I��/�<΃ٜ�8{���"�[j�y~�b���"/\Q��#3�=������/l��(-�����ݯ�����SZ�/��kPUH���+�"�������i ,g����b��&�5i�'͑�j��n&��"�1|(
5��7$[hr���C
�a[��0�B����=�'r�?�6��8-�#ϙ јWHq<�dA�(�_f�J҉�X	�������vj+?�iH�������pl
,�B�����&�ܡ�.��g�1grD��~�b�%d�qb=�5*]��/ȸ��q�p�b�o�C�p"��1ͣi �wƿ��y����ѹ��M!���z�� �|n�#���h�%�l(���a��Q�@<`o��R�s?j�h+ф�=06Gz>>��<���� �Hv9�I��S�+d���%�A�N��-H��1�-u�P�{�H&��P�N �"pw
�Q[Mec�z����`����vxL���r�d'֙N�Ϟ�Ge<�|��z+�x�Té��_��ǲ.̶V��==��t3tX}H�@NBL{�u��J�pK�oM&�����V����}�~�����r���BFH��S��p��h�#N�%�"u��='%ƀ��Ҳ�\������f����aj�O�c�c��&gN���eFQ�I�k��M�a�ͳ*�l���/t@����k��XZ�����D����<*��%P��n���I�y�=�UA氪�U E�R�Jb��9���s��5Hڶ��Fz,5�ua����ȝ�VW��Oc��� ��! �O�$#9��|�@}��Ye~��Ģ�]_�4�?�D%_��W��"b �w$�6a	D���	�*�[��$�'����!�!'.>aIʟB2�Z��T�;���h頻�'��쥧�c'^.i�1w�e��80�V����qjY��맂�cV��������I;{�n�nj�Lˍ�$U��6#<�6��o����m�Ț���)8�"�lY�"�8"����1Ͼ�8qfpZ�~+��;脂�Y��HG�pQO�����>�)�0�Di/�OGt�P���Ϯ��(��:�YK��-�	$.d��Լ5P�O0K��`���Ň'[��%fqIAB�~�����O�<��*��ʸ��r�sVO�j�f|C����)p�_6QUǅ=��g-+өG�M�� �+�BC�੿;<�G> �����Q�r�EMy�_����۠�!F�������zr�*e�Eo��&���E�  A���m�_�'�OX���)��_��1�K%�8@�Y��#D�8(�&�&	)5�0���h�-'FoAx%��
{���*����D�aދ�(��Y�o��|��
"�1\�W�3�ݲY݁�'V�<4d�d�r�|\�<�a�1P�'S�0�Ջ�Bs ����&ݘ���2�%)��W6��v��U�Rq&7Y�����
$���R�(G%�)�x��M��w��T�3���H?ض��U�
�Ӻ��@.�ɉ�G7�o���})� >��9�!e\#n�;��ѱ��}�@T����n���Ns\�!C�Kh� ���WP��}�cO��Jϙ��o@�=�P�8+� �Ն����p�����&�|��M	�M�n��B}��2�o&E����`' 6�A��l��?c Q�2�\ap�dG*��4���='�?�(6�
#���,��-NmHhl=�Ku,��'��Z����
�RI�6��|E
�n�S�~� ����?Glor��-It{��36$��|�}�~�׎n���(����� '��EN�
��
HNd�8Z��W�̠vA�M���m �=3��_���yF�z8NN��H@L��I�F�p<k�VT�"�l� ���t�
SY�"@���7�VJ/���T��,�a�w"S7�a��E�s��
���	7Ha\T����X"2��{�UQ�U�-�z�k#�B6�ȓ�6a�G:Ni�q5m�N /��#n�i�5�U'$í�+Q��lt:�zD�5�bRA��WxE$��j[m��1�2{ uDԌێ�X��w��]l���/��,v!��d#n9KVo�	:�"�jl7^����J����C_a�ͫ�Uzt�<���I`a��x�>���LE��Jr�.{Ƿ�>�5��˫�=�Z?�?&�$-��5���e/����K~<��|>%I�U(R�w�s	��wX�'N]��o�֔��~|�m�����_4/a�OE�9Rx2�(�,Hׇ`1אa�A��j▨��.v	w�;��<IjO�7��5p��
0޴ɇ�(�������*(��&�q�����>}n�`݀�D��r�뭐����m��d�E��6��P�y}��U��a��`Q<Q���|��&
�J>��u������*8\�s@�xuLDW�ҭo;�?��]�rvW��C����J��H�By�Ƌ����W�����~����O���� \$��}���VU���
̊`���N�u]>�1v�)Q艖�ܘ]|9�o>��WqN�ǐ��ܑ�-x%��Sr�v��Zdc�gOeUTOn$��w��%BCP��zZ�"�B�埧��v�����t֘�W�>ɭo˔�3�b@�v������e%������^�BZ`�M�k�#=/�]�k��6�$����m����E2��"7 ����)B���2�=a����ˌ���c4K��*��䜍Z3��#����j��O��*�;N�? (3˞u=�����1*�Y'#/�J��naǰ��L���x {U�W
7�QCb4R��zL�rCb����A?_�Ƅf���whLDa˕�T�C� B�NW��L0k���Fv�=o���"�6Y���XM���MF��=~9$+���^i{Qe#��`� q~��)W�Dh�.BRte|�d�[�3��9�\�l��`ɠ�c�o�9���ײ4��;%5wj}��7�񅛼/}Qf�n/���Q�2��MC7̌�Ddkx#c���H�_Iq��"�<;�bz���nX��j?�ޞ+V�5md�VZ,
��p��=|��z1�9t�QMwf�
U�։J��D]���c?j��~+%��
���`9G)N-���+��Xr��2%�����s�v3.���n�A��Ruʭ��s��!TR�  �>�}�+���*ZGzP���jkCqa�.&�i�B���򡧤B�c~��?rE� ��R��~��S�\�֛1���ؾ^�g�Қ�fv���G��r�:C:8�|��F�����_�9ג�c�~E�/tҕ��{�+M���4�����\Y�a���{��y�B���t��9Ք&6)��(:>^�-'4pxg5s�Z�9����[�.2�[�KH�a�\�cH��l�{NW��R��"琬�E����u �r�N���r:58�<�4- ��b�2����O��o>��g����1�q,XBrZFuW&��$y�tM.�3$j)Kuw�2��[���E��������%��`6�z���"h센�@�̹*R#a_���Q����SR�s=�ﰔ��]�4��Eq(�����O���b{���*������N�ʹ������l�wގj�~Ŧ�DO6#p��&(���Lu���,<�����-�G?,�gɐ�z�?����ؖ��0�wƪ�N�Zp�O�܀-�H��.��IU��%�3�O޴�q �{�����%���6��HK�?�7��O1~��ߤ��ڑD�$D�_�.�y�I�L��PS�?��X�� P9{e_�m���m;�F�my"b���p���4u����
@H���PB3��6[
��_;���4v��Qb!�z#����%�Ь��!6�r��>M+��~�G]��T�,n��Lh(��pZ/�/>G3,�;�V�vgm�ҭ�6��'��z���5�`췱K��u$RpG��cUѝ����}� cq�:])D;1����p����j1*"�U�	��:N�،��Fx�zd'ؾ�e�!�8#i��6&�o]4�{%�8> �{�F*W���[���˙U0I��e��J!��CLn ��*B�'d�b=-V��ĭzFz̢��{2]�Q�� �����uĩ��d�+�ߞ�6��C(z�׋��e}ak�+�%��Cׂ9^k��|����C�v�^zV5Y�)�1��U�:��}��6<	sr>Aq�hL'$I[kIo�ך���]��>���:Xַ����u�?������o�0N��2�i; ����hN���m���a�Cs>h��0N?sz*W�ot�rZ�D����W��cV������~-k|�~�6��G%S��N��ʶ�c~���r�w%⛂v��.��ò�WW��Y��B��HJ@�R���y�<t��V4��Gb5�s�ThsY����Q�F�(��h��K�_������ZE�D<s�JYlK�?T<�;�Bd���QO��c�t��w���\R���Q��lL������#Y����X�_S��D$��M�jk����`��@�H�Snz��uA�79O���|4H)�iޞ��y���\b青xЕ�K'|4�W�0�yw����y�˙�ǌ�\�[Ҳ�|d �߾�\�u�&��KDm��Uz��FF(E��s�LB`Pm�%w'9ŷ�W���F4�(vR[X�R"���H5m��_.*e��u��t����Yh��`M���k�7�Xq׈��ʃ����B�e�����C�|�g!>'��K��!��sA�_L�dt�Ss�0P&�5 !��a�A}Krp<2�dY.�[y�J�׎�C��l�U�y��h��qf���0$��o��s;o���D�τ�a�=�\E'��� k��-�^�� ��8U�=�-5������}2U�[�Q�R�Q�d��?�4tבR�L���8;���r���N�˶o2���s�o̹e����r"�se��`MA�}	�)�؇I���l��>���0�jg�f�֓38�B*�Y�9��"�RݗǾ�# ����>�����;fhe*g�:��l~���E�5@5&�0��
A�u���6{v~0V�)sM	r�29�� ZF;B��R(�(��q5��ȸ�Z�4�g��D�����,��d�]q3�Q����/���pR�+���`�kCUh�,6�2�W��"D�&�}��\\�p��g�(v�bHc����8��G���5�E�vJռkw����a"�5����9k��>K��s?y��2]� t9�;�*Dd/���2V�t�G9�]A�"/Νm*?c�쵆;��w��b�� ��T����##W��$��;�k\��ݿ��_��҆祜��ov,���`�r[XI�o[�I���i����(���@�a?"/"��mɍ�~|Oူ^� K�����s~3�6�w���XL���W��C��)�o
�	�V�:?�lDroP�ՠ���ҧ��o��'�ż�>�)PZ�h�� �ݚ!���=�Y9�7R^�s�=yYK8<�v{��3�&�7Q#�n���ݻ��6ȸ��j�9�݃�H�����^�@['��>�jažư�gU��� �ܰq�ؖ����ׂ1t�e�)���5L	��k��hh�Ik�:�-JP��C�(�An_J
1�I�7�&Ch.J��
�[c��H�M;b0��p��P���^��d5�J�ܮBJ{�_'��r`���bEl�ԕ�a���X� o�O\���.�ގy�%��e���|RȫPJ��ж
�V�oף��Z�VZIJY��bߌ xͯ�[��~��ӕ�g�& \������9��)˝�����F��&��;=�ܩ�4��Kߨ�����4-'0�)h6��Í�9�Ŷ8�1�X+�<��u��ȼ[�G��y{�%� �Y]�*��qZX��Y��^��X��>�A�b��R�p��1��&�}y�2~TI�%�wT��m=�+6��N.�������"�$rq�v�J�֏A���4��Y'.3�4+�K�}�}�gy�i���ӱ�Ǯ�L��0�+�,+Lk��pG����O$�Z<u���d��Y8�dp'w��^�jdG��ܱX~���N#�(�,�����lc00���Ɣ.b���� %d4��yK*ځ����?�sҨ�_*�������$M��׏����W�.;�\��2�5p�E�:�$�J�=.�`<�Ί�r_��w�j4m���BS-:���i�r!�.*OS](7[��\e����� "Y�Dbǽ�X%�t��s{���ǿ6}��?��!k.�ߐs,�
�x��=5��D�6��ހU�&u��aY����i�zB�]����r����]�mR���l{��;��}YX?���8WGq��9��`�:��?n�M�x��LƆ1G�q'Y��Q���l,�Ս�����G��2FL��^- - V���s�L���,��Zl)�̣�rar,� �\/u��Y���OL����9������Q�h2H��1�F{��N�n}:P�^{4�k���މD1�~��;]���a�dK�p��\�zr�f�I�F�F��nQVT�J� T����S��:#�+�|�]�.G��F=1x��Q�����=�kK@�tS.������o�M���6���E�I���ހ���+ʾ�b�ס6֚+��^Y5�wci��YX4��r�q��M\"#�MNE�p�{$\[w�>�^^Ue�v�����@�ԚBnW�3��#���=��)��ޘ��f��K��u ��;|�YS�j�|A�_q�v�/���=�X���f�u����j�J��d�(ާ{�'�-{6yM�nfE����O�x����
-b��b.��7����t�7��#{�]�]xC�.��<cUOD���k:s�����2�>'1����2�>a��ua��n��J�FwS��!@��Ug�VN�z	��5JQ��w�G��,6��D,����mx�c��r�[ZVX���q�z����Q�\����tKs?��1s��o}!�w���(�+.HB�X�0ư�H�'�"\��a�W��~	����{ת�W�fWCTZ!��DZ�*n��ȵE��<F�|̭a�f1r�1-���&�N3�c<nm�,�z:[3x���;����y�5&May�o`�I���z�H/��IR�KEI�#M�\@ϣ/���d�e6V�u�B2��hez�w� T�b̲�2���p����GC�$���g�#(,l{�����JZ��gr���M/�ji�Z�H' �&�VH|������6�滋��
��b ����p������g�m�-��R�8%�%��r �,  d*9��Ǩ���oqJ���u�������D:ͥ*'(5UM}(�z֕�4���Bf`�Q��4�[ZE�D�ħ��:Tt�����,��8������߽#�7r9����Y�M%ɮ��5�d;�/���.�w./����7���F���gZ?�J�v/�-T��W3Ћ{H:����T�_�+��w(Q�4�:��t�ҟ���A_���O.�H��"���Y��E�I��
��F)[��]E�����Za"���@Z��+,��u�|H����H�*ߧ���#���M�%h�y�����R�H�D�p���>a.*�k%����5i�	D$
a�q~�pK��ے��7���g��s4�`�� U��R��Y�Wa�AsjFN�[��d������2�y�C��<��eY�Ӆ�?����,�&e��V#��F,�<K� o_&����Ž�>r�����k�w��Z0���ȃ��<η��
V���������TU�F�=����FrN�a~���l�oR9��v7�S�M�X��A֡~&Q��i��E��=�K���jV�2�b6C%��>��� 7�"ȝ]� ���n������dVMw�uDG�hR���;�j��T���s�
�����>h�r�`٤8��_�d%"�%��5�1I'�|��gd{�=��^�K��ñ�)dV�~�R�0O�����C9�����q���ԑb�0�|R|v�4s��a�y�q�q�ӑ`�,v�ZV?�,j�DU��\n�����P��I��A}�|R��⴯=\��5���6TW�{e���� .����E�"(iD�
�\�	�j"	�ρ�M#ma��=�F�/0�.¥o���b�Hp��P]�� ��5N��ǦO�����C�#��iH���g����w�'f`<��
�-�Á���z�+�fg�Q���x�jV��@�k��O�G�v��Č�.�"����9�Y���� k�RS[`�$H�s,�{3�� ;3b5�K�n�c��51���u�j���'�S�,�©�g��zrn�u�fF)��`���@f���'����\��k/����k�2��Qg��L;6
����γ��R��t�Q�QQ��Y�*�����=�7K�k^�Pz��{piY��ƴ������8��ϥ�<���Khȕz��Ѻ~��=��\��fT ���>咱�EfdJf���J� ޡ�u6B�Q��&�}���D@p�#6Ͼ��Hz^ꏲ.`9���CAF-�/� ��~ƚ> ��(fȹ��
�; 败�Z� ����֩����\!x!�+��M�O���"��p�����lk�r���|���5r�<TVDx�> 
c!�T`"�,��R7$Y�Qx(�1?A��M"�h	,>g� CZ�V�Bx��˩E����F�	:�׫A������	��T	���@Dsd�\�6�����\S�ѰʸD�Wz� q"��C�o��a�v��k�W��Do��	_H�Ə��b{;N#�B�q�}H�U}F��и4dSF+����o?���/ڷѣ4)���D�,�)ȵ��T�!@<�"^����Ҟ"݅�[9w�2cWz���L�����`I&�ur�T�/G	|6�2J3d�BH~�i/�TrH�s��Om��o:"!vӑW��O%�!}1�R������&8|t��9�����al�x�C�����$+��5T6�'\37 3Z|��&��b@;w�ʌ��'��;��h�v)�H���V�s��c�bk���� b&�s&1�ōT���x�%����7��T��Yi8ĵx�Q,�^IS~��F�hXG6DE� �������V��t{�Oȕ9:ʐ�V������'��➊�D��h�E���7q�	Y��~�&͔��g/R�\4!�m���п���m���c����?�p4L���Dl�A���9�	pJ��WVñ;����Eھ��,q�&�c��Ġ����Q|&�q��?���w��u��3r�t�-�+ϣ.�۫����mOѸ\���f]\��1�|�|HC���y��~�ʆk��w�v[�����_Ӎ�ma؀��[ԛ�z�R˴v��<&�i��C��-��'�K5�#+�t!�c[��'�H3�;+K�6�3:S>�X5�a����(˄צÿ����C~�L <�_;��8�Oi��5��Y�Z.�l#���3�@V�P7�
ԇ�o0t2'�i-I�}B.�f֔/�����t�2���E�B>��2�{���Slm��/��%<���y�uD�V2,�F�	5�ǋ�5���#�.Q�L�x>���8�s���vy5@!���(�	rI9
��Խ$��h �ѨI�a�h	X;M&c�r~lF�; ����Au��8Z�;[��q{��Wh-j��K�Ā�bwM��#�.e,ѐ_�'d&�������ܶ���E����
`]n���O�`3W_��9wS�Mkrr}k��<MpJX`
�M����*���o��L�%4r�~�i�g�5��7@��"�UzW�@�
^{�ϒ��Wz��B�[�H��aW�j�~�����A��l���[�Mn�����pz�;���Ǵ�b�}#������V6Pl� �%r�۽)����*�1$O<>/��m�d����̂+� g���jy�黜��ě�}(<]p �o�,���j��qNu���AW��5Q��nwv}(�Em��a���ٻ:W���p�JT얙�M�rZ�)���ڛ�����D���E�["�!���i���k�%��J	\�&O�NU	q�T�������eXI����� /6���j����sƝ\F'>�������bUE괚0|!e>���
���э/�z�����QҀ��ƶ&;�[��-s���+@�/��U��`��DX!��j��]�;N��6;Gpy�9�,�9�;sv�,K����+�W��.8��zr:���i���ߍ�$"*�O�w̆���s�%�clg9!�]��Ҏ9�V
�Q�tr����l�Ueyi��O[0�tH�L�5�^|�)$�oRcq ��=K�{(J���n]0�ta䦌�܀cde���#��k-U�с�'k�,Ͱ/�D�E���Ё���#�3#�!}{ �JF�|*�.X�>8J��d��w�9i��a%&ֆ0����-Lņ���"C�S�:�$���eҕK�����B��x��nZ��ܩq�G��!�y}��	\1D�ɩ��TGnP"S)�Q����΁T�uڃĤ����eD�{_bц�\���K��bp.#�s5Oq��6��32��}G��g�/0	�q�o�� ���򍞩 v��7�tG�c�J#y#l�La��{C����~P^�!�����#���|3�T��Q��rd�	�3A�OcBJvh��a�A��t�@g�җ^��FD��؞�@�=z�����ִ���%:�E|v�\�|7�:� ]G˖��^��t�\��o����T)8�cF&q8�k��]\��M���/�L��~���z#�-��'��P�z���4��3Rȋ=�2Ꙅ*X��']��J,4�O5�8��R$=�������h�m��q�d�p�wמ�il�yxc �4�CqAg~�nj�Nd�m9wJM���{v�{�z4���]�Ь@�8F���#(8dZA�YA���d�z ;��ף����~��(��z񋹸���T�.��+.!�/�q�F�P/p��V�I���dD�)��`�L�8Ѩa,�]�CkX����M =�0у'EѢpĕ��å���g?�P�Եd×B����묶��h�5큟�hV@��n�6�ޡ6�Pq�]�m����z(�S/�4����$	��pT޶�{:h,�ҽzC�����|��y2�Mm�e�����\	Wrb_/5Ꝕ���8���a}���]���%^���6_��8M)nIA���-�l�a���P�pϓ�	!�rIǼV=K�N���]:&���6W̋\�zx:�8��w;�(I�	h�M����?�����|�7�����k�a����1��^��I"�b���~���Z����т��]o�}�M��iw=���]sM�1�g@JP����*t�� �4��ҵ�ߚ$��]��Mo�����4�+��h�fЂX+Y�;��0�+�iܲ����Π�@Hm�]����D0V���4Q�$k^��(?�!`>�dT������gh�nkUr�@���3��ֺ��O�U����&��E����@���# ��W��� ����CPJ^P��*��� �&(��V������Tz I4d]����׳��`
}�̻X"����?��qt�l8�8��8��ϛ�٩�LO��� ���{�Fl�b��ÒN����g��{st(
����8�_����ԋO5&^ ����p����<�sOܮ�[�L�`����M�p�Vg-���Κ�S��?A�%�����c�����T3�N}���t��[�Ch��ܐ��zC@��mB�#�rӱ",�^�ey�$0dvn����MQ�~7�U�>�J�����5&��Ml)=�K_?�^�ӿ�p�t~�BH;;J9/&FTD�p��D!2H�����!x� ���66����ƫ����(�>�c�9_,�ή|�xe��i��g�B	a�,��Wf6�.bd�g ;�_���0�u�𮄌�Ӵ�ӤUO�Z ��_3���+�<,��=r��g��J���X\�叆fK[�������.�A�O�2Rd�T��5
����Z=_Q.�ǐ/����ܦn�����K^,��}vC������=��4��ё)ckj�Pq����-f:�4��]�6���Ζ�׆e�d�r�2�V�
m&���H0�o�~/s�b��K2�������Pi����4�Q)l˓�a�2/ļy�,�oaM����y�<�N�ހ[���_��^���i��ﭫ�WF��˖NC_����)�oo��,��{��Y"���D���_��������}�� q`��L����w�֨�o�.4�o���s̾��[�)]99�)�v��V���&��A��j��3��X�A=�TB;H�;��l������+��DfI��U@FKo�?t|�J�R71�sق�x;5�=`�8�ȶ��Ồ�)�72/6d�_/%Ā�k��;���n��an2�1��#�D��z���K~�6I��P�����vP��B�C���r��=�HP��o���o�g�^��eB���a����Z��*M;D����䱂߫�D���5��}�cU"9JS���"�7���i��E��m�ͽu�H�� C1bܱe�{��'��FvUЖ�KP��+����`��`*s�� msM�γ�� �̚u�7�5��Mkc�E����pϰl�ގUJ�7*F�O�*��2�3�y}W���U�L�/����셤d���&e��Y%~?�̿�D���V�h��Z!gO�u@����v%�����E��[%8+-7��d[�� KC��}#�y�i�R�� ��e�6R\�	���)�Q�L3TY�йd��ڨ[�>���݄ΠxEO&Hy%�i��ue@����n�W9Z$����%��bL����E����p�;��;�E��e"#i:��*=���b`y&؅	�+WǄ���̈�Bf�E��!d%e������⤢N�g�&^B�pf�5���������A��Jߕ��Q����y���x��:�y�嶌��\d�s��H�~dR�=���qX�\}�1wP3�G��?B[�������`*w��r'�([b5X�K�q50�~nk���v��#�3�ܩ߿	��D?ا��m�UU�zh�$8�z��gm��>��
G���X`���ॹ�zzu�����v8F�'m{�jN�̽`	F@�������rX(8^lx���g ��h�����V|�Z� �����	{��� !�������a�-^jm�4����u	_�P�}=i}��@�4i�c��G��k�a�	��m����)��Y�^T�f��\]sZ��m<���+�_�Ԃ�<"7O��R��G�����"��Uk���%*����*G\�X��z�Ģߞ���I���%�q����=���ZB8��f�J���؁����V��ei��3u쑰���Zt[;�D��hە.'�����T�̱d��sAଅ���A*����'���1��|�����Do4Ҏ��i��7�溵+ka��[�n��!<���O���*Y�pECG	������3�צ)'y�ߊ8�5��J��{o�Is�ۗ�N�,�3��? [ M�1����Yɗ	��sZ�ǩ\�]������T�DSw�~�������*<ۊ`�/��"�$��\����{�A�%N��N�����b�8�J8�YgO�o�C810�XtNn!��-I'��ȟ��6oPu���9���~!��H���E�P�n}��?�^5���,�u}�w9�e� ,f=�
���5�L�7j�;]�5�����;hK�%w� <5>��	�4��h����~"�x�&?�B&As/P��DV	��[	��YEmϝ�+��؛��9 D��]>U2�M��	���π�t��	���C��G�J�<� d�t���l�����zΐ(R��{#óyvM�H�����M�1Դ}k�(ˏ�ͮg�����e���;�Ss�O �0�y0�^��ߊ'���#��҆�?ߟ�ǻS��m$9f�f�"�֒��DM`>AqV�o��x�;�W)'�������0C� ���NFo:3@�)�c��^��YtA�8�}�&����]V�"0h<mw�]kק��*�U�)�G;��U�D���zɫ2���ʶ���_9���U?'C!��z�L�b��өH�1JVhrq�^oc*����f(,�y�Ն�u�x������0�����0�%*�w����X��/���f����ɮ�����F|*ּ6D�����X<�`�$�
,����g���a������������8K������*C���N�͸x�ʏy�9���v�Lq�+���=�;�Go傖�a��ުmq!'�R��ݷVOZ8��d/B$;(4<9�%R~:�WT`����K�v(���u2�@�_1����3����I����"y���`������}�W�:�#�y���xa���Cx���dD�&r�D�.`��4v-�"�f��y���3f��a�R8��\��Q"'�f�c��
�5k��Jw������L(C	�fKs\QD����/*���,��fxp.��qZ��WJNvtSES�㚗@�iSB���(�p~m7����S���7 ��6 kzFiZN�:�[q�*��h���i��eo˵ۤ���V��U��K�����,�C��S����Q�l�� �Ƴ��W㪥�t���BpDeS���o�Ƕl��-��#ϰ�c�"���AhV�zx�S"��$��\��Iי�i?�q�ǵy��ۛ���Y��`�>�Ҋ��F�ᡧ-{y2U�&XM�'~����N���q�K�8@��ݦ*���T�^d)Մ���$�����}��U<�;��8Ws-}U�)}���im�V�T��\β;7m�4�b��5����~�q#�,�`&)3��m�1�"6��^o(2J��(.-;ӛ�Lu�֢����aK��r������s1�t
d�� q�/�*Ha����n��஑��<���H�8L������Rn�gW���ttlr�s��aEB�~�+֐��T�r����Xs����8X�3��j#{����nI��[R+V�]HK��i�����G�zz�_S�gtyv�D��e�\�b`��f:%Bu�R,x��dyAB�.����J��/ ��wǏ�$��y8�怳_�յ��h_�M;�@��B�{�?�&�ڮN�ɃFReTT� Ž�����L��1���ei�~0<u$nA�����������$A.��UF&Q;AD�d�b�G��@i���4�����r���:�0r�"�K�N&ڮ<����6�,�3�o�4{��ƶ�1��D�,�g-d
��[���y�u^���䊡�RH�˃Mms[���X�f�tz�P�iՁѠ#Ԯ���T�n[�7Ĳp��t�7=R���Q�	�]+�_s�IUb6v���0��D��-�Q^C�lF��I}Ri23���+0}�fSԄ/��B�>I���s������@�.l�	�KxR�gF$/���@"�.�HX��m���� UM8#��|7�ȯm����.' �+��/j�~�`6���=���AxY��v/f���yy}���&�����O�ɻRV�'���}��Xn�d�~qUw*j���>���}�>h�7��^�2�`0w߾I2ۓP��
��6�@�ߨ-
D���v�b�/�լ�6ۙc&�0��[���h�!5H뀲V)t�D���$]:�}��A�8���tOC�V�3���SQ��0v2�ڗ�ԅ$���6��[
�Kse�)@�(\��K�������d~��8�(|ɘ�)������$��d8��H�9�O���e���6���B��M*d�Ӫ������4���?���5)��#/�V~m��Z�VS��ݚv��8�yu'�Ư�f�Pǹ�o�l���Ύ'���
����/K�bZ��OU(���~)�����e�����19u�������﫪����2ҐG-�B�	��n��)�d�=�;�I�"F��T�6�ލv7���<)#��ϲx��FZ�s��e�͑qs�[�<P�5G@􏊎� �%jBe�U�n7*!���fb�SI9��|�H�a�.��MLS^��Lٲ��`H�Ty�;H�@�Wkbe&��'6wo�7��]��vɿ����b8�Ċl��_&C�^Aq�����IN%O ��g�T����=}���lX�L$o`�m��~*A�z�6c{���3j}L&e�f>��fZ���������C��y�j�"Ol�j����,���D��&�'����j�̪&�yٳSN^r
?�֕ '}���"ZE]X��ǨѴ���g��E�8�F5p���w�؜69�d_�Pse[�1�aDcG/�DU�W��#NvQ���X���r��]���=�U9��Y�|����s�������<���e�6{�(��ӻ+.)�j}M��)_:��n�[�˂z߹v(�-17c��^�e[��/��Em�+C��D�(&Ƥ��IfQ��卐�#�)�j�A�*]���I&vQ�6��D��01'|�k��#?}�:��@?�g�D��3-.a�x��<n�\I@�'�0�����*�4m�z�Ν�-̣���T�����ؤ��Ů�H�˪��dm ��1
QP�v�j��m����z\N|$υ`{#%�7]E���J�����e��S��U`F$�����L=��*�z�7�j�;s�v�K�����?����2���T<�{cʯ2{�$�h�;����ܔ�>�������>�&�����<��\?'���s ���f{�	�uh�J^6R��9 g��7ztIv!�����\@=�L>P� �B*tt����ŀt+��⟯�e�
��8(}?.~���6C�:2��}�xN~��ud�G7l'�[��*�2���|�+UF����r.}D[�4#�Y���%�f��bCi��;�'J�2�q�����	vj��c@X��\t2x�@���;� �/�/��b���9��lP@���e7S&�g5��J��� ���q j.7��r�fc�� -�_DY��$���v��.�3Ed�&�qє�t:��@<tEf�_���
#�g�~��N�j{���<)dFGu�ziqo>$Ԝ��jI<��|��QŞiOY���~�̍�3�6�N�
�U�5�U�
K����ԙ�'8SX��f���Ʊ�g���QȘ7���Ӷ��O�ז��&��y������0EQ���w�fK��]D��܍hz�hmW����1W��ݣ�����r����>�9�2�o!�������F����U���Fܒ����	��~+�/Z�x哨�ʌ�&�Q�V�&,���|�z	+�y7n��|v
V�́��yp�Տ�K<1ЫW�$j݇�1|-�2��)Dhvp).:��g���l?W��V܌�x��ڶ�97h&�v�!��c�oJ6���g��,0 gMr}r��O���_^�|�3|�1���0l3�v��J�z���樲�+m�0x��[& H��;
�[`�$sg�����l�z�{6�>]�N>�z�b��˫\��\��2cV��������?�ډ�jZ5
�Mp���V�5[�&��i����݋Ti^�*�,#PIx���ô�ܒ$�T)�Rf�'^5vC��ɪ���ۻ?�&Ԩ����2��_`Ns����2�,ß��́��'N���H�\�MT?Y�]����5�0��ԋ��<�|�����	"��O�� ��S�ʎ(*��X�^��Qݏ茎���٩kp)��=Hm�|4DJӘ9l2�,졻�����蝤�����!
@��9qތ�?fbC	{�1h������j������� j9ưBbD���Rq��ٲZi� \����No9����g�#]U�`X���\��>���hdM�ZOヅ����K�Y��	�8m'_����s�!뼛��YF�.X�a��c0�=��K����΢�7�m�v��А�~`����|�J?�D���֌��&�m�D��j��O���9��8�/�g��)0��yrl����d�n�$�d���G��<"v��.`㒯�q $A�����Ǜ���O��<J��\�.+���)�f�I�p*X�6�W|�W��6�Z��<mї��iA}��/�P�b�#Ӎ3��Dt_�.��ǕS�!x����r9�pRυ}�y/;�ѩ���j��#F���lzը���>�*pʢ��NYé埻]W�j=�)���g#H�'.���AR!#*4v���!� �L��1B�9Ma�p��
/���W-����iJ�b\�fz����$BQ;D�\���2� �G$c5�;-��qe*��L�V[/�\_Vܚ�%�(ck&�S�%2��t�޷�t{�UE�qL~�=�d�|��[�wjF7���	V5����z���po�p�'�:F��:0w]5y6g��M�{	��~90c_-d��1ET(>lT�:#t��'��.�g!�����1����{폽�NF�ȯ���/���_��(�s#}Z�&[�i�j�y:����:̗T0�xO����W3��Sbe	O\�o�0��!c�=�
3,�����%  %�!�����+Ӛy܌o�o�d�������>f��g���-�������`g%(���}��{(��N�p�]��Z�_,@F�n(4������r����h
t$��;�09�\�F}�Ѷ0�>}��4E��쏛胕�;rTp�����i��i��t����!B�J,��p��L�G� @i*��:���t�u���z;L
���f:H���|�vs?��k�(N�S�,�J���W��"5�Q�Ѻb�b���3�\a	j3s��!�Zel]j�x)�ռ�|ϤB�?TYT���qk���$����ᫀl@��ws�s��U!�i���$3��zT�*���)�%��Ne?i�}ɆI���n�n���!�i](*�At�3*{��TctSƐi������S�ɣͽ�ӳ�o�Ϧ-�]M�0+Z�V��y�JU���|(\
ϝz��.���~og�����d=�m;!8������c
��%��n�ؤB8�:5��r�l�_�kռV:{�S��n�� nl����{�Z���|�P�P���tV�h�mU9P���4��
�q�n����`CT�4���N�0$eq���O�Au�K���3����qn[��C��+!׏zqD�;�u����3@��ȓ�xE��-ב�H���c���Լg{���1���%~���yH���1A��+�@�U�كű��|��e�R�-�H%��.+������Z�uo���,��gd�4`���1�e
"
��fG�X���M\L���5���ϗ�}�����z��'��X	��W<�#�q+��u`�;��Z��Bu<$c���;���\�1u��5��L" ��̎o�� v|>���,8 ty�k ��W�L�X$���|�U�����΄��М&�}y��2p�Y�{��t��'';�9<�K ��f�
`�l0���Y�q����6�?m#�aв�!e{��+�6�{�$D��[1���?ƨn���fεo��qk��hZ.s'��q���?�f����t*�?'Ħ}��n-��<<�ٸ���������<��O��Ӭ)V�s��Ԋ���@O�HZv�R�����W�_�1�������:�<bx��#��0+%ݬ�LT_�ǰP��M��M��CZ��[5p��B
��<`��Ԏ�u�C�NZ3L����]�\��S4纐B?��O�ѽy6�1���,:���*>�Hk=�����1�t{M���N-��]�S�L6X�^�F�I���>�EMM�n���4�3�$�
<���z.�����7�HR���[q�z ��F�;,��^1a�U�Y�ɳ$,�t��4���iWqq�������{p6��3�ߏ댇��~_��uX��wt�C+_f�)!y���^��g5�K�� ��z��*�80�
Q��Y�a�fl�`�a���k^J}ڹt'E@HX�J�zc�w�wѷ�a���rSO�������rǤOۤ	0䎖�s� R9������!kf��5v���ich�&��7�M�y� <{���!O���D~~�UM����Ƞ����+�W�[����Q(�u���Ab��i\���� � I�Ԋ�l$3)���)����q�$���v�BƁ��]�#n��|Z-Xބd�g	s��o����3O��P���v]<���i$=��iq��vG�ԭ��"�jۦ_��QYS���лQ��C)��O�yk�8�"T���p��/��ML$n���s3�KL)*C�V�������+0)TFgX�v/��Y�Y2zr��< �+��·Eg=k�iF�_@��7VXX`*�/0����"�%vެ�u��-^���诖4*|�����N�33X���ȗ{T4f8�팻���m�ڂ�C]>$��P�1�f����Zc���%�(�;��	}���y)2�JΙ�T�xs��\��A�H4�E;�\3�:ޘ�0�Pj�G�|���xK�Z+�X�aQ)m��wwn��rz���WL`U#>'�k�Lx;K�rXF��u�]� {��=�1B�/q�c�У��c��L8ϲ�y�̰)7�d��/F1]��Z�4�:�.�����qjݽ�M�����6�A܀!����>�=�KM�#�ɇ�8H��0�br�vi+�;*<~d��/2Z"��Q����ZC�j�Ú���2`��A��,�a���l�bE��~'~Ko'��b��k�Ծ ��:��b0R(}�6��C��K֫��1(�~��G��լj�PFf`�#D�ަd͋�=�<�Ȱ�o��<U�&h���_b��08}fGv���쉬G�T%
����Ǌ����q
��N��� (9	Z~��<�N��o)ݫe�c
re��H�������Sfs��P/C��d���<�X���0���'��w'��DML_�.�dfE�*�Fe���%-M2���=`V��&�R�F�_�l�����G>U��*�򓒔Q�@K�5��z�9� ��lgEV1��.;��ata�vV�Fug��iR�'�Z��ooB3�Zѹ����ZW $�c�'�~��8�,$���L����m��)\�R<紅���L�+0K�����o��z���bZ=�I&h7n�7r�p�  �	VیK�G��޺���>�n)	�w�����/�,��7���m�EJ��B�0�BT�G�ƮEU��z�¥p��'i�����W�U*����g�43j]��]���]uv�ą���_#2���6V�5���챔�`.<���#�~�U���7O��M�p��6�u'ggP����b����GT�D���$h�L��߾���7�a���d���&T�� J� S��� �����C}���&,X�` ��Ki� e-4��k8����À�I�~�s����<����1�&}���D.��3y�vG�0����!�����oD�dnb�#J��y�=V{�%u�f>�����V�F��WG��K2,���������cp�5T�@��_��fvUO�Lߌ����ŷr�8�I���Q���h��&�p���(��JI�ha�Y5�t�T��S��W����v��o�$����U�5M�Q�6����n���	��2�Ƅ���Ly��*'�z�������f�ʚ��
!f�%�"f����W���Nf��Ԫ��/s7�.���e[�^����9i��PY��I"7�/a�b�c^������%��
�5>����z���'a����N�r����=����r��!j��\^}�e���š��xj���m�:3�K��M4`��M��DY��GV�
�#*r�h�����r�f������u�Z-���Q{����?#��	Ҍ�u����$F+u,�p?��	.��v҉J�=��H,�qp�	� �C�#����U�`b%T�%
�h���Ϣ`�$_��D�t��g�"m^�ڙj��|�{v+��
��,���j��IA{��=��M�a��,i�-��ؐ�k�m���L6�ܻ��"����+$~�]`��=*������mL�4l�J��pӺ�0PP�,���Sky΅��R�M
���K��1�R>}�&J�� 4�f�Q�������U%~�*|?YjI'���?����f(�ml�r����A����~��~��qN�H<%z�(1)Θk;{v֚D6dF��Qf�Qɬ��U���r������ե���~}ЕEWi�q�;��.���u.�iv����3))���uK�7ܟ���q�u��!�3��^x�-�&my��^�����JuZ�d[��Lj�`5PA�K�܏�d�U�ya�K�}k�SaAm:4L� �[|.����%�Y��R8�����ʡ�2�9��$�rր6;�c攱M1�B%a�]�==��暎�Ûz�\N	pk���Y�{��a���]#Pe)?�!祮��ʉ�w�RP���߹��
L�)J[g�\	%F"�wP�x���jH�0*�qJ�t�;�q^�:�g���a?+�9#�,���(��������xw���0�'i7$=���J59`8��BwA�܄Z��l�b��g��ť�ڶm�b*�,<(t�$-�M�>�{R���բ����������؍~���hy�9?��9
ϋvj��e��^�[$���'�o����ҷ�K=|<V%!�>p�1�����zS����/YA��	�
I��RxY�E�y~��F6�Y|�;���2�h�O6�Y����g��?�F!6M��9��/5�Y���E���-��{�!�7�K���M�V���i��r���C�&�.�k��N��
�xH1����'�DP�SnEi�����Qb���*<X!R�%Oxdb72=U�D�`wgx�Kǖ��x�<��E0<�3�AJV��b�/�=�S�p[9t�tA�g�!%�?��%_RZ�{'��y�*�٘�W4�G�DZ-����2Nh��2�yV�T0quM��f���v�@s��VA��;�R�]!d�-�ҥS#��/�B�x��>����+,ک��ߑ��O��X���(n��� �7�pi�
X�;j���� �����۪���pu���&((�	MG��G�^^�����d�L�'�[yN���Ww�F�u-o-V ��3���ⷤ�*��Z�p�+߭G5�Sa��OS)���Y��0y�A�^(7��Y���(���]��	<`��d���J���Y�6�DM��5hp0�N~}�͝��\�%W�,7��mg�	)yAs��WԹ��@6ܝ�NJ�nM7P�pOJ����k�$;i��@F�wڟ��S��m��ϲ�6��SkH8�����J��E`ɀ,ˬm�(~�o��b<��+�X�|�]�Uɱ����"����(�p�����H��MV�[J�%�5H�=_�TP:r��|��%�jd̉�T���sL�Tg��\Wb���;	�_���U ��_
��k�T�T���m�$\&���b>���w�,�ʓ�@��h�RU�~T�`��\PɼM�ܧ�d
���KG%���J��k2��B��?ը4�#MZ�cWK
�k#*����[���b4x�[���5���NQ)�-ީ�����K,vcǜ�x Nm�o�kDy���nm����O��l(E=;�)8�����LK5L�r�k�?����7�U��Ȑ�r�T[��6��,#z����ep�[fQ���|?�ό��{�[_, ��g;�MGq�b��ukzᖂH8�<�|�vx�������7�S��j�.4��2⎝YO���HԈ��K�J�0A���(փQ6k%ߔ-�<ʟ�����oP���DX�>��u�$g��Wz@���,����Jj|W�I�K�]��-���k�=�s>c���A��˞Ͷ#W[��oZ��E�U�`]uK\E-|᠋�O1�=��Ǐ�Ʉ��=��i��{5�R�5�(�aR�lU����/P�1����c>5*(��39]s�����I����
�����l�,V��>�W��~��9�RV��A��ǣ��a�@?[d���ȫS";��v�����,�ʩR%�WD&c"�ݛb�O�,bu2�0;��4%�E��#��l��r���f0����-�S��a��M�d� _u�P���N_=���2$��A�ǭ��<i4���$mC4�����a}�@�1� T��'�|����� ��	-Q`�P�[tW9����ؕ�T��Z!�HUQ�݇����/����Cs#qԬ"�V0ؗ$Kǚ�:iU�[fP3y{�2�!�%!;cD��%�9���萲���ڍH�q(��3���$�6ϛ�[Wr�*Gq��>q�e�(�B��Ow���|"��ХB%]��G��	�M�*�i'E�kP�g]�������Ũ��f���B��gF��Ί�/����x��iz�Ӱ�<�=i�ehp��Z�������Xc�%`)�"V�BCVLA

)��!=�"X���/ߕ����s{��������k 0�-�"�
қ���+�h�ȸ�B���w7�ya�#%�Ә��^�F��S�/?���s��ϊ��ǀ`�ћ��W�O�ETɕ�b�JF_��g���_
�"Q�2�DԇF���e�6�ͱ���S���8�~
�κ�Ќ�j��e��Sj�>�D�I��?��#�D+�w|e��B����̃�y��K�5��-�j����?�U�2]��n`���#�X���A��)�r����Ͱd&z��3��^�̣�采<)iu���S��}czEjw�V���nl�N�H��6�مdYg��J���nME�=)�s�M�UN^w���g��Q�J��6A^���r=xk��
���'�d�ʚ}�x�3O�lFw��!����ͱ�`��C�NfF���4��N�u�"pa`T�p�1$H,�4Hf��A>�ܝ�2-_��*U���ǂ���M#QI}�a��m���;��?J��p�lOo~���Ȟ_ovbWg�K\Y�ZQa�S��DM,c���6|�$�W�n�Y�����*�(�.�8{�tf[Z�>���b�:ʿ��� 񸄥h���v$=�蔒o���z��w�O���6m�;�1<I�0�:$Q��S�+��l�	,^]U��QT��W'�D'j���}�� ��C��\/ғ-\�����`^Q#�>�@�4�K�9���ؘ�|�#z�nb��d��[7�х3�pZ����;�-��n�2�.�C��J+md��J��0�:r�^���b���IQ{���a\�dl��%F�K�~_�G3���p�1!�k��7������E
�iZP�� �-�l�GFh��̲F��B��0��A��P�ڛP�]_��rc�qȗ�蕳9��o+f<��p���i�����d�aB�yl�4(>^��76�l�S�&A��b��C���^8��=lvqx�������~p���ܺ#<��;�rG�ϹF{Ny�ጃ��@�;2`�1ѷ �	�{$��L��Np#H�I�7^7xڡw!�so�$ ���Y���A��u�Y��l ��A�3>��֛�}	�'Zm�k�n,��Q��µY���\�� \����fНpz�'��kܛ+�V'�zx�Y>�	��,r�#�������^w��E�<%��]Q#\^8K�M�� ){b&�k/Q����d�\):m���F �u;���$L8����E~d��� WNa���}��3Y���>E�$U~aY��'~��rl��׈g
��6Ib�#�\Zo{@��p�'=y���������z�q@�X#�&��C�alӸnv_�k�~5����Q����[�v�[B������l�,_��d�(�i�*kZ'ȼ�P�(��	���-[�=/=f���`��x��E����P^D��m�����])�z	����K�~8��K?ɗv ���$I����},J�d���y)�JKY#��&T ��B�f��V��	l�O$�K!�i.��X�m��F���Ś��� ����_�`m�"_}�gw{C8�P�-Hӹ��r#j�zu�#�y��m�R���:�RS3�	wI~izjyMw�-~G� bw�7M� ���u�'�KV��*�W��}"�훛�h����Rʧo�Ut� s_D� �FWh�u*�|��vY;��Y�_�L5Ed0YMW޽Է�v�;���&��U�0|�'s�CZ�ӷb�+��ګ0�N,"a�﫛V��W,+��Z�b�����\Txާ���{�_V�0�X��i��gFaø�m��)���H�(O��慍���t�hЍث7�ΩX�Nf0�}��{U�S��O� =ٲ&A%�a%xF�gU5$�h�"��;A�`ߴˑE�q�l�у���|#���`��#�)\�v���n�';5
.��a���(�ʈ��ZO:�h���)`���s�,��3*^'^�߃i��͞�Fw��ľ���;��V�{����E��H�%"�{�ܒf���U0(�D\��ٴ�PS^�6���m-�6�:DUp�c�9<f��@���� ]�,��W#�;ZƓ? �؞������*����V�ş��͐
wJ�Ɍ���{'<�y��T�q�{�M��l��i��0%q,I��E�����a��w��u�����R�D��!z6Q{�V�ݎ\��-����L&��v����3U�,���j��-5���3�����ew��_7�k]�^Un�b��>J	��$)�ǿ�0���2�W�<\�[$����z�~��\R�N׏?$8+��'C⾿Eԙ�-=�Mb=;+��`��`�#)E�S;���4�s��V�}�AƱ�6��1Pb�-��?]֔�h��E��,� ����n��������3���߰���XM`�YI|7�o�����h������+�x_�^�q��}R,�����_�pb2�	s�w���4$u]��bCX^�Q��T�y�X��}.p*�o�,�9�.��_
{�oK�R���n#���乳�W1\X~��X����%ܗ%�J8���n�>�1I�`��k���"A��&�N��.9=�9�F�@4ӝ���ԅyB�:EjFetByD˪���8�pj4���ܳM�0	���N�-�;tP�z>1cT������� ��~3�,����I��&Ad�0��GϞ�A 6�F������ʟb��_��M�w0�lģ��ב[d�2 ��)��`�K��^��GU�y?H��S��=��b<A��fS&��Ɗ�������Nt�@�Ro���9S$a);Oq���]DЗ��$K�Z�3F*�ȶ&�1~��z,�e�]2��P֮��e'0p@�_����i��>��
�z>+�z���2����yhV��^ܪY��+�;(ܽ&u�*\��#y�#qn_�ѵ7Y�;k���h�U�����؃$��K������	��#0c��Ǝ�s�?�� /�zhE<lvMQ�_�ٱ�/��X�Ԑג<��?y]a��Ww�ȆԸ���c�*=�����k�P:�?���E2*m���Ǜ:CQ���|��v�yթ����anes��G�  ���j�y�s�hIco�\>"��"�J�R�G�(� �8�`b��l}Dk�W<� �ʐ�O��C�W����С�;�)G`�+�������'@�	Zx�M��:�0�#���f��� ao��E�+N�t�����Z1��II	���>r�\UVq�a���\w�^�$�&='O���z�iF�  	q?A��IQ����U���rJb�T�z!z.���r֮��m��0��p���]�:F�M���̶u���W�,ɔ45���X�����8�W/D2tg�����G�dn�Հ���v<q4$8P�����V�W.�.�����[ݛ\chOR���OS�F�� �Ԍm-�1��49�2���B65N��*�ړ�={�����7�vb��Z¹��K��z��9EYCY�$��p�a�>�?�u�J�E�fR��>=Z��t�`�S�P�2 �W�gσ6��B4�����|�[���S*{eW�I(-�Y��d�֊!���K��Zd;�7����&h ̃'����L�	7��pN��ht]��嗭����)w_��.�1rQ��� �sj
�e0�C��%ړ��3�h 2s�{@6�n�r����w-�����3���Θ�g���`w��n�R�����A/��hr�l3(У1-p0��(�ۈ��uW_1�
�f����խl����`��Q�
�C����(�M)�Y�

B�?��x��l�@��*�?x�PW����+�;�20Վ����S���҇,��a� +��2��l�aSc�1�yZ��ó����Y���{�CA�r:m�S�֖D�46���C�S[������d�Q�����a��
��3v� �1Ƶ�*�ŐFZ��ֆ���K���D|~vܯ�o�0�:v��֑���4�_��E6�N�ʦ��{@�U~q4T��UK�!Ş	�A5���k�rׇ%WZ�G���v�Ɯ~��Q�q�8���_��GF��<C�?�|Iu�I�oIc_H��x�JDd?��"Y;��gE��<U_Q#e)����X+'-�Q�h=���w&@�EUĠ/E��ErI�P��.����ܷn���}�V"�gZ��R6��[hq5��*�h[�!�A�
�s�1򲷪�G0n����}��p�m�YQ��B��vb)��u]D-b�W��>�G�O���pp��)b����4�w���ɋS��Ѐ��E0VoS&n��-�RU��M:k��:pnq-G�Q�	��r�٨�'�C SUG��%����\�Q���*�w��h����v�K�����4����]��ȡL��V^���@#����w 4n��O�ׂXޱ-℡�|ޙ�f�1�TG�7&y�����huy�,�-)�W����z�H��m���qGzNǯ�eI�V�.�����J$��W�a� �,`�U���Js� �Ʒh��/m�<fk��l6Ϻ��c/��Po�_�M/.y��gW�?~��{G/�k�z,$"(�v�+T� $8�;k�DH��oN��m�}��y�s?�#�4�]7�K�G��c��V�(j�{��"ɅZ���c�Cs6�G�/~��OV��U��~PC��IzTL���\���n4��B��v�0cQ+��6��9;�.�ZVۦ���8#�c�!�ut�*���;:"c:k6�C�8C��3�z���`��L�u$@�攵>��M����eC�[w���9Q����>�x���lS�J��v�c�&Ɔy�18�H@��+�U�a���77S��׌x:��<����r˗ͫ����;�����7�63�'£? ���߷j(��z[�p���*�C�D$r��E�9]�G�~;�#J��=ZB���3��~�¥^�33���?�k�����n("�m'@�A�I����[�q\��3�,��e��߄�m���9�β�[��i�g��u� ���~�Y�\(7SӬr,M;�>n�j��$��|	�K���)Y�J����u��HPIiA�ӛP0�����cЂ�Ԝz������7�z/�,ο6M�b0ۛ ���=�!��3"�8���C�u��ᅧmi��j�}�-1E������D�U�M$�����=�Eنi����1�]D	�Cr�jf��A���CHR��Z�h�MU�9��l�Z(쪑4�3��83��aR
�v�.)�����u�v(�;����{j�;���Sdr���F�MoyM:���\KՆ������/�`O�PZ8&+�T�s���M�\N�t�z�M�C���/�l�ػV˾�2��%�µS̺�ۘ�/��}�
���K�iT��<���p�%����=`Ƅ�V��/�Z�C��a"1�jEﶲɰ��Ne�p��)��*\�S����hL�Y�0�9����e�k�^�<�aT����ږ��o#���_ȋ�+�/�^���0���HZ-!-Ά��Puk��KG/�3���B�DG��'Av����>��`�n�M�Ä�4�+��5\DAA�BH��P���ȱ�3g���B����8C5���ףydO��a��.dLPꮇ<��Y�L����o�
�颯��ADc�<>E]���A$��ڭ"~���L���:땫>T ��є���ƴx�x�*��.�`4@�\S
�\' BkU��mz����mi���8��y4TFu�z�kdV���c�N��-H����zGyu���DЎ���A"�S�əi/q�������@�s1��Q^�3��jo39G�3�xB��&P�u�~Y��~��A��1���^��6���M��Qz��Y����S�������~�#z�=�%��E[��O6��|�N����B�/8y�~��m��2�z={3�����,=�~S�E���o
����[�]�_!Y���*;����ܔ����F�5�G@��-�;����� Ό�X �$0c:�<�Ѿ�|s�fnxS͍�0��� ��)���P@��n���\7�-�����A�|j: ��n���/J2+��(�����K<�W���)V7�z�в����Y�T/��n
N�9ڛn�}���K��(�h���Kqd�����7�?�͵k�_���!���0��m��rҿͭ#w���!���m�v���e�i����@��e~�e.�]�i�%�ȳ%F�H��5�TfM��/��S����2S�D�P5�BXH`:�:�����J�5gW�Qc�lv=\ic�ݴ;�y$���,��vƢ�ViR�}��OY��E��5�B����W_Hp�s�s��]ۧ�j�<{=�[K���#qs����3��7J��[��,���F%��?�۩�b�fh����pO[��ڿ`��`��Ȝ�QU�����e�A�n'Uv���N��kP�2B��س*x; R������"K���p`Qɧ��0	�J߳�N^k|��N8 �G@d�Q#DQ�HL� 3���ow�Պ�|�]z��7�8|%��L�sv����j�Rc�iN���c�]!cZ
��
>����.J��锽�i_c:P�gՔ������;d���^���ތ��M�L���#��o$|OŅ��H�~L��x98W8S2I)i�i5���-���������j�J��".Y�y��*J�o.�(��:85�*xsȷ��Q�V��<4���4��m���+�q���.�RO�fUw����	����v5�<J��b��/~�f�2�!1���K��w_1����֖7����^����l!�z���/7��ɖ!ɷù�3�3��#wto��=� �Z��l��:�+�t�����'����T��)ƀ�b���|n�l"��x@���Aւ�ׇg��3�:�1@Y j:�Z/���"h�W�1)�J�����M�'���	��(n-p���J�X�u�J�Ⴟ8��{��I�]x�RJǇ˳����X�O�� �I��W;�㩮s+>��g��S��6�,�̭>&C�\�l����W>�2̻E�f���F�y�{ffR{g�s�I0���G�nqg+y�q|$��CW�T�۶�=����!��p�v�lw�k��j��>Zt�t#��l�?�$<��˂�����]��;k�qP4�.F��E�z�+v�&e��}O1����ފ��!=�IS�R�<��\�KD�O#����|��+��=�š8�Υg��J%��i/ad�@U���]�&�$^��1i��O�[��2�j ��iܟRW��vA�⒪���g��&����D�u�`s�o36M�{J�,r���!@�����/��|�$.a�g0H������V�1`����c)� �w�[Q���C�qU�^�B r��o怜\��v��`\7o���I�ށ"��E����q��&��C���Z:c0�����i��k���<�B�r�P��������|��p������L���W6�x9�1���0�!��%8�H��t�eT���8}+t@o@u�J"�����Er������
*��n�4	L�1@�c��px���������6|1[3T�m0��?�k���q��/�L��Ps�8w�jy��N��m�'��+���6�����w�&	2�K\�)S}Fրv�F�IIR���Z/��d;o���q/F�/��X�ߨ�c�����C�/�@��e�	�,��)�0�M�*O���'� ��DM�k��V�]c�����5u_?�[2J&�TLc�t��`[w�;����` k�i��u�����'POd��Sx��ZU�������:3V��^o4E�v�f-7 at�"@�h7�]�ܤ@�E;:���H��F��K鋎(w<뙳�T�X˖��e�`�M-��w�NWT����$��#���<�l�_�´�����BS�!���o7W�:�+�r�J��҄��Er�`vL�!��"ɦS�ܽ��m���a�@�a�스�OPU�ckG#<ڗg��n��-�E��l������OO���i������Ҏ�&������ǿ#���U��&��x��`\`C����>����%�+�����Z�V7�gY�;�AH�7b��5a����_>�f��5���bյ�&�(7=2�~����"ί����bG�^��Ԙ$M�DU�@�J ���Um+�ȭP��;!��oS��U��[��S��H�0�j�$�������5-�L ���KY�e�'P>�qjl-��o9L.EA2�z�N���!�)?��R}�:���f.Wk1H��F�3��j����b�ޕ���y[�űĬm��:�r��=��$�&�~'$�sF�L�x/�>�[�/d��b�<c5��0�b�3���� ���!=���r(/q:U|d��u�K�0����:GlU�QI�`_}�ϐt��!i%�za�ُaLz��*Q�kf�wq2�r[�v��ĺx��w�n�>=Yh��`<!��{\p�6�x�8J�%]������=Y��F}���\m7��޲Ӓ���e��vB6�ps�ցE2�z�g34g	�˪6J
���Y�(M۴yH����&tkh3~De���؜]~i$��/�}���#�7�Ľ�e[���~;Q���S%�Iyy��{�i@NT0
�:�2����� �󤱀1��Ξ������9c��24�cb#o�;8��/�x��JLQ����P5�-[�:Ao7���^9Y�]�x�	]ǓY>p).t3f���s��k2�ǽ������vR �΁�����@$�
G�k'[�5'�#�����q�"�Q�,��.;]G��R)�QZ��Au�q��q1P����c��7Eq�Zb����C��U�bt�"�A�����[���x)�C���Y� ��/r�;$<����@���s�8�����_��	�����'�s�@�Â�}u�ظ��*ˣA��^�n�F�@��:D�N���\���M���­��ݼ�l�$�2�ĘIC�k)����IZo�%���wE�l�u��M��k��!�޳�3!�'|��9u@��;���f�����T�H���X�tN�OgR`�w��_���xS0�k/ʄMm2a.,�+`ԍ
�����\�N�'u�,8����Þ4���Z�@��|c�z~����kg$�Ƕ���'yFK���׮	�l��Թ<������<0
p��,�[P'�=����B���<E#Zy���:T*\�Q}ƹ���it�tr����rGpY.��+���h�h�		9�v�s�"�y�ŉ��S���xQ���l��������Z��Q?c2ĸ��W�=��	^��Ga�p����(�61��§ y�7cj e3�"+;�.�����S��'z�����̀b� �����p7�B!��?4�ÿy3š��V� ��<Nm�>
uS�t�-�,2U6�3����d��
A��:�r�|GÑV�NY���� q�Ύ��b�'"դu�	:x��2`���BI~��������>Dq宂
�d�u�S�,Vf��t�-��zkd�*�-7���¨���Gs*�떀�u���xD�V ;����C����������\�%ޯ=2��sC�r.�YǢ�g�"�1èmrP�F;�cRy��"�ǚe���z�ˬ��;��H׮����M��_'-��m�O
�|�=Շ^F�4��a_Q����^�����r˻R,���ֿoC��~-:����WJ�-ZM�=B���翷�ak�p�Z��J��(Xʨ��m��# i=��R��j�������H��5��΢"f�|=���T.����-�����ɽS��La���U�9P*���&��Y�|�v3ڟ�/�%�Ӊ�)ocu��
�G-5Z������=T��IUΗxY�4v�O�-5�.�������[�2��������Q=��g��v�g<B~��X�ũ[�@�V$�1o�5̄�EL|��/k���$���;��0�`c��ְKO`�Pj�_�U��9%3p�ʠ���Wꪛ"	F�F�E]~���̕Y�W-��yk]H暔ކ�̒���N��τ���;��0��4��g��g���8������:M�{t�A�@e����郶>�a-�Lt=e�y�� ��}��#D��רP���HЈ�n��FZ�:��Ԩ��Q����́Ӥ����H:p�d|�C�Z@���0�	��v�0ܢ�Ҿ�lB��@� �Y�^E���M�F>l­J�"�[�����[��h���)phK�yD�Xv5Z�^R��;=��@+*]w ��AAO�������g�`8Rn�S����Jz]Ɉ'*�uZ���7X�"V� �N4V�:�*�RHxkNV��Q��J�L7�;� ?�8����d[�b*,"��=��c��n�5*e%%\����f����/����
"F�:
E+ӣ��g�jcl:� ��l��6��S�WKe�ҏ���4�|S���\X�Z���4������ �FMY�7��e�M�_��$��qa-`�QT��h�O��.�F��l7P��_��9b��̴BT��Þ����zʦ% ��z%�����Z �l�����#�&� �f��<�-�&�͘�9.6~dͶ*ׇ����p��Z�L�b9��gz{h]�|&�[�uȺ�%�]f��`M�?(v�g� ��f������b�X
�I��R/�_߯ �)���f͔춭���x�i�N<�H����a�Qh��Pz�Ů���0�/3{A%����8p��9^��z���.�Z��V�6���(���v����B�U8�~���8�8�͕����nd�|�����{��%����fz<�RH�H��nrT��)�¢�I
����b��5���
���5�I�x�1�Y\z�v�J��(��;-����"�>�vrk@'����[��Y`\�`XX���V�R���/�Y�$�e��O���K��,y��G�#ٲ���TF�6�%~�6����άV�p��_�{� ���*�W�0i�7`:�q���~��]J��W�'�h�ӵ]>4����,�3۵�$���Cf���,b88�'O�}$��w���]��ʐ�}7�¢K���ؕ��k�K<�YG�熜�CP"S���[�o��0d<֏,�A�!��^���T�G�M� $<<U[,��8��jVѕ1;S�[��;{L��I����A��z�"~|\�vo^������73˔F[|o �<��ɫ��=�������C��<+�J�z�ؿ ��`�k�g3�<� ���em���S߷"����Nģ0�0��6��u��DdZS� B �h߀�ݔ�k5�|�}&�Ö���X!pFN�5�,F�yZ�w}�(=������Oc��KJx����L����Y�/}4ʣ�!��?Y�� ��n��>.Zۤ:G���e��K��� W]�i�]]����3-�ۅ�;
�%xĲv���l�>�V��aI@�%xl����]�znK{-�<�8e �/�}M��`NS�F(1E&"�]Yd���mt�"��V����ނ�Z��.-�9�L*y��%Z���%Z�"��~g�N�ю��q��O��5�:��x�'}�d��wSX��J����G0]�Kk�v_�
�bC�2�-%�-��Q�6F� %ٵ�n�Tm�	(�ea���s\l��S���
X�;j'��8�r|��xKJ�V�B�_���n�u!Y+4y~��T�v��h��|l*,3�Z�x�V��cO��_d�mA+�W� +�MdZ|9�ݺ(�p�	�g3�V�k� pjS��A�o�BrA�Q�~Q��� �eRSb�l06,�?  + H�w���Ǎ2-X��w���v\F���0�Ǳk�����M�V���������F�s�z�����q�Zs�CT�~h�)��ݼ࣊�
T�l���`�4H]���]G�T��#�a-����0�Y�;:�l�г�v�2��b$M��^�R��a�#���J�r�G!�7�w�90�ߕ��]��'.@�eCm�e����z��n� ���edO��t�Ќ��ꙷkp�|����{��m�q59IȖ��},��:<i��0�G����o%���\���;0V���lJpCdu��������)�/R' a�|i��.�^̶�ܩH�g_F������N�8��l���� <��	s+
��]��enU�^��<cA	�Kw��«l�( �0���r�.���)۷1��	Ty������rcΠ@��)5!����Q�����C�i���M�^z~���"M�yڛX�,i����}G�EH�<h4�f�)	��%��"�<�0�[���d^��Z�s��ϣ�扚�2� �x�Q��I�oZ׏_�aָq�|���if��B?��gR�Gz���&<�Y�D�8\7"�MQh0*`�	�W0V�ۦ��Jg�`����n� �$�[*�c���z�yD�]��S�)�E�0źGp��y�L��}�Ԡ�Ģ�r^�?��l�h+?�O��1��ǟ���4[��
��2&?̸}����A}l��O�y$������+�?&v�	�U
T��J�o�{`5F*�|��!�:("���B��WZ�)�|�bäR���29e@�bP�h=���곸D�@�4n�ao�������d����:z�j�<hR~|�9Y*��>y�50-oz�z�!S��'��Q̉�UwP�,�ǟҞ�cLr7I��k��`���Zse]Uy���9���Pᆳo ��T+�t)���;�5��8����H��#�d^�Zx�x�s�Fv��t*�lQ)�Tx_`�s��Z&��`P==V�j?��jio�a_��t�Yf�!�M24�l�"@͑]V���%����_.������,o�xn.Ig�� �@	C�����z(��%5	kEo��"��ÿ��-i�J��a�'[�V3�co�����u���܇B���9�97lA
̓=] ~z]@�����v��^[pz>�o0��ڒz�Lώu��� Im
wg-�J��(d�@����v���6.���4$�6�������"� ���:�	�\��\i'gW�JK[���g�#���*}}���R���w�`�C���m�s�غ�Z��t�`����+@� (��VGĂN����	��K��K^�U�E�nk�� 7Z'��C�h����8��f�%Hl͠���a�Q�E�TuK �O�WÜ<B�%q���Oֲ��uk���Ï��?�˗h���Rr=~? c3�f_�҄��3v����tT���U�7~��� �'�x�U�����qw8O��)�m��K�)��SO���"�^�����1Y9�X{��:��K'���J~�# ��7!OT��;5�M��b9�1��N�T�ҩ���nz�A����p�x�)�^���׃�c�KG"��`/�/����V��[�P�l0���K��R81p�����BH�b۠�)i�#j���n�wD�獔�IaR(&I�e-^7|a��\]S�-BZa�3���-2p�8��H|S?n�юt�
�K_)*h����8f���@�;�\�즐C�{<+�#摔P�ql������t++� ���CT�L5zj�"��}@(MpR��8^[*��}t���8�y.� YZ5�Y*H��w��n�-䒈BM�
�(��u��r�<[����$�OVa�!��[8�E@Vw��4��S8*����>�|?�=TT]QarRMN4RO�A��Qq�,�ݵuA�vj�)P��\1�����Ri
�	�)�<ތ@[�5�Ф4�U%F�"�ǧV�4�0��E������W���$`�]<|��BVu�ƚ�Ɓ^d�M����i�eWCs���@��tč�/��X�&�4Ÿ��"��`��j
�A�G��Ǵ��1�������:��,Q ��}�
+�|�vX@^�=Z�{��'�ޤd�0,Md���4����C�d �鳍�Y)��eSU�>���$�Pvb�R�'���02_�̗�M���ĻMY,6�<���-a$�Ɛ:<�N�O�HT����T�����3���\Gk�a)O¯��[���xi#���r�w5����l~"0����Z� ^�{l��=� Y{����V,�^@p�V}MP�5;ugSJ��'�����c/$r��8�pz����(��A�I�z0�7��_�-;=�P��'��-��c���GW��~��e!�^$��M:��)��_{���e���[�@��'C�I�Dy\B=���R]���GA��Y�b��@�=�����Ѕ��5��Zf�i���Z���;�L�s�x�ܫ�Lʽ�hVy�������b,���ړ6���-Xl�I���Dy}��u
��D�Q�}�洡�d��בN��0ћ�����OY)8ٕ��Ԯ.��8J{�����[l�7}d��x �Ϸ̥F�G��n�,�G�mh�6(.n�F��W��;�8��
�L��؆��x�����F~��b���K�c� ���!*����TҦ(�h��O�˃B�%:�鹎��N>E�f)��	OvzN�V'��>��㇞�W�Y�f��k��K��- U6���f� F����jP�����I��$�y"���!?�D�ҥ
����5NKӚ�Р�i/��O��s�+�N~Ůcmh����ȥ��(`��*��6'qi�.�!@"����.�?J�%O���W�����2��r'���?4Y|����Q<R�U{m0���r����XJ�x�*�����߬0�t
�� Di]щ7?A��ep�Z*dXᅇ�7*Bd<��b��JS&2�~|��"�[oHd}"�����/x�v����k%�˻=�0�`�=ٻ݊���վм��жo�tb�y��� $u ~= s2��:�>�=`4�H�w}�~�i��@�5�]���|S(�5�c����������g"t������y��J��!�'%��V�
r�ək+��`�<<�����o�@_���r�Se���#<C:^ ���k�Q��6���inI$��%����bq���pP|'������v��T�f(Bx���aqrl�o�?9Ѥǌ�Ǟ�)
s����^ڪ����(��I�~���nAh�h	B1�q_�5�P,��^=��'G�i��[j�K�V)CE�٬���g?���B���|��t��M�c�;{D2q��%4u7dm`��WZ�*��$޳�<�kuB.J�)�ү����`arx��y_At(-�����s�>�mI�V��+\��4��|�~�\Qת-98��������]�v�U��r��o)��:���B�D��,T�U���2����́�F��tEh����<���*�!�TuXQ�!�o��W�V&�?�&�s�Mb(��L5��Lg���mc���J(�	�ދ޺�uo;ʔfY�4�`�fg�st��7#;�����Etƌ:x6��va��P��-�i�|�T�z��DbPj^2L���������M��@�S��`E�u|�Yb{��֡&��
����%����U���y�lr�O�u!�&�7%~UX��B�k��a�ֆh1o:�,z2�{Ӻ�<���Ao�K}HJ��\�&��E-���X\W 	� Z��*'(s;�շ�F������M�c���m�n�P'��'u�@:�������&��,/�ϛK8~%���/�0�s��_� �]��� y_y2r�`�n���m�o>�<�]$�̑U�s�+�U��w��1)�\c?u���&�9��k�����!�,N��q�6�\�3���!���xg;��aD4�z����:$���!�tPˢ���#�k�^�dd�U�>�_R���6[��Ϗ��F#���V�o1�i�5��h��Í�
�ы/�b�A��nb��=\%�V�{ٟ���-^ј�\�]�x
����x���GY�G�(?���@�!�L��)s��֗�m�n��=
�|=��6*��2��2�8	r_x�E*����u�3�A��Q	O����WV^�isI ����,�+�UG�b���������ش/��
�d益?���1�8�� x%^���ܱ݊�=k
��3��b�Zo���F��4tݔ�%	�S��PN�_H���)�+-\,�f�c1��Ƽ�\d	F����g�!M�
uё�x�1�������L1�������CQd�Qۊb�L�f���)$/�q�*f�)��y�5%"�ң�j��9��-�/ݵ����TfE�Vܐ��}�Px����&h�BG���Np��b�4Ot�#��9L2SX�����I��Ǔ���W��^�Z���w�i�)���Rڟ=4
�h���N��X$H�f��$�
����ۂC�d�n|f�q�%ߎEQ��W78@ $�h�V�b�g�� �l�B�v�BRi����P������V,GE��K���τ|I4�8���F�hA�M-q�5Eb�A�q�������:!�Z��t����˞z�ڜA�`���dM/�ʿ���k�
Ə��DBCS\��sT>B�-u�:�%��[�4- C�w	5�N��W�6����2Q�-��6��V��Q퐒J��5$�^z�4�����������V���-(�!H�Y��
�2�s�s&h��������M!���)���H��n�>���q���S�K�	7�׻𵨍w��߱�����@d �V���}��P ��z䤰�G��KL�><�z�o�;��^;��
h�+��J�S}w��=ܛ���g1M ���ì��a�`:�������C�8����^n��a����&�S1j���9�A��y��
���!�C�75�c�?5B�p)�Z�4[8�FK�{�L)��s�$b���<���ҥ�|s�ݖG�!|�!1��~t4�$��=l$���/*�$���	շ�Wz8�2�c���nA2R�J��
�ķЬk��MN1�OҋV,Ll��s�xў�"�{%�����Kw����S�k,t��ʟ�s��x �m3�M��`�I�-(��ͽG�u%q�^���p�N'�,%?�놗����H׸�ǟ8�}�F��d�7qz�|qϙ`F���#-����>�C�Q�Gޅh�N*{.K��[�o������wN�������������~�����Hޙ�Q���Z�;��9˷|��3̈́*1?w��<�:�N8���c����"֒�s=ʅ7�r�VW�n�c	���b%f�� !��!H�����s��r�}B��r���7�s8RF�1oΖP�L��6�uW�Q�o���7�.IP��w֩0m���nv{��8}%����_�n�f������zxNR {�7�FD�b��7��I�I����X�ǀwq.<�[����0ϙt���R�#�%ߠ�����k<��.�<���٩�/�F�J
.Ro
��oV��RN���z�(~���v���<L�)	<g@�O�ç�Q�ٗ�j�X`J�H���=�����p>p�@���H�Wf.��LNGz����!p;�!�Nْ��t3���'.'����T��鷬mW�/��������n�UJ9��Y�d��x�D�L�cpc(�=��>�R��l/zi�s�O,!V�ǂ��x��<�"����џ�=rc\���I�Z�!�Γ|I���)F�:�����5۾��u#��E��g��ޣŔ�d���L=�נ'	��8��RR�.N!����F�L�{����ϫ!D)��m[� �jo�����+-��/2r��s�`�G�M�t�Ɨ0��4J�7�at��փ����a�,�[�%��L� ��Q��0�\����QīE4L6Zg���8�*��0'�0"��;=D�t�C�`���x��KO�&���\O�3ݹ�����X��GG� �sf=��y.z ��k�q{J��ܣN9��ҖeS��ev-�3:�%z|����-$#��0`��9�N��(��ܪM�8��p ;�.�R�?z���u�5�5Y�,��!���a�j��eK��[�$O-ǂ���9�g�FC���3��äj>(��lȫ��ױF��j����=����v�ZI��3� ���r⅗)�)���-�T]�
�񱗀�0�d�������[�D��@kڪ��B��e�p^G�=��e�h�ý
��
���^�k�y:�o�t�B��C(���E�ѠV�n��`]�$q���a�ʾ�O�%��"r^������X^�q(�p8Oˋ�g�f�D| �?q�-�����<F�t�>�F��/���H{��6�2��b�Ѕ�T�i�jH�XD�;���&��Jp�����Ս��m�3'����1*Te�FR��?y�����#~3�M�+?
"�G'}��nM�n"7��߰O6��r3v#����nl���u��d���<���j��R,���d3a.��k05P^�9#w_Ñ&�My��F��'҈��v���]�\
�H�.�K���k�V.�"�{�^�&���2`Afz?J�����v�o9����� �u~�(�]�@�3T6V,��8g�� �R'����O+mܼa�z�(�����e�e��8�Nm^��?EQri��t6���������e���� �]%?~D�WG,���J�X�B�����_��M-�ނ����)]`�3'(g�k$����5,��.��j�VpT�_�TK���F52\���aQ��7=�h�Y�o4�|ʟl������%���ƍÏ��J�2��rH���{��_?';o�h�h�
o�e��|��ԇ����C�I��=�L;p��ǫ��aM&u���S2��K�"(g��d[HteY�
���ʝg_]k 0Q�Qix$�j�w�b�{|6���2 3Ӊ^TY��͆%Qt���fWWY���jPMnE�k��`��;��M�q̜k�i�S��"�?�������6��G�%����h����|:�Bf�ܜ��3���(>rX~�NV3���j��N�$Iz�f��|t��f���%^>r?ν�tΏu ��A[��mn���h�[��ϋ0oX����G�%��r�i	�u����Wl<�Ŕ%�-(��1��3�x35K?�����p'��6�;�E(9������������VW/�SN�!��B�bJ��w�:�m�E�c�qj�ܕ�� �2ԬL�*������%���FC����o����T/%V�yϻ�O"qk���x�F^��E�YJ���rp�#0�R�n4f���b�F]D�tԧ���N�`z��lɕ�>>ra�hl��t�^k��Ђg�m��W���J3�7Aq�0�1����kZJ�p��g.Z�꛼i�M%U<"�cj�S~ 6\�q�t�M:v���!(��EG�C����0�D��B׵��F�}��]�,Q�㔴Ƹ�A��{�qcV��X֍�7y�i�<��~:!T�<�j��!<8���Pij��bd����{�~�k@X�A�м�C���oM ��4j��%\�NJ��*����Z@�/�w��B�\�>.�aK�>B(�S��sd������GS�n+n:p������M��6��r8�հ|.Z yعyi״:�]�.��\$_����Ü����"a$	���!֪I�X �����ٳd6�Y9�}]���PN?g�]Tf/�j%0Q�z'3'��nW�/�5o�|�
�u��>8|�3�¶\ISƬe��,N7�/�YvY2ٯ���uzS{WnL�b2SO��$
���#~�F}�i@$!��$o:�0%�O�H��,�"�}�	��hB�_����^]�����Z�IԐ��b�yԷ���)GqBkf�n�-��4�����!Y߿�3;�fr^%[w�9�n�k��V:��#ƷH�7l4�@�nG�g��D;E��N5j��<����١!�c</7��/��'DI�����6�������Z��T遜<U�E�μ�gf8H^I��M��� 3Ww���&@�SB� �ܦ�J疽�`�.����b�ՁK'�*dً���Ѯ�q_�6Y�*Ƞ�w�z�M٦�6�jXފK�Dn�
�H:�M�ƃ5ǟ؍a����&�0��7�o�~�@<�h����R��{��>�i�}���<����f�[�9+�DA#�@�1Viq�sMC�raBhD��պ�V��������K�=;�I�WTS��Vz�8��kMFKJ�=i��@Vț?���\���ٱ����^�����שdW��QF�����룀;��P�Z�򋈰���)�I���2u����i����wwZ�A�0�Ŝ�uق���W��}w�E�5���zE�M0��ڶ��ݳ���r����A�8�Ɉ��2P9iNK�8ܢ����5'Q�*��Yt[RU�g�p_t�M����4ь!�3�b-#������"�<NL���33p�蘊ςz��I$�{ݒJ�ۍy�\VSp	��$�q��D����(��Uwc�p�u_P��T�E48,�����9�Q*���.����uw�X���Y� ����s�!`1�n;)<�=>%^�ف�oۥ��4�J�1|C�!v֎�$0
���N��a8�0{�T`�;w�<��W*\��{)	���(�7B�^
&�*ò�1r5��#�q��F���:��	ʳ���Y�?�=ץ_2	����U�RY
�R�B���m�]lZ �:�8�����>&~�m8εij�h>��f�Y^�V6rݫ����/s�l9�A�]�.��h�9�Z���Y�)2���jO��M� �:|"ar�f\"f�;���ay���jg$Uh&|��Q?*�+v�����_]?ŭ���'���<y��ۺ�b']RGv�(��r#I"0+h೵��3�\F�j����GEIJ�;U�گG0�j�����X��:�
���*�c�?O��I�c�N��e�o���Im��D��@|Bk�E}�Ѫ��X��"p?F$*�w,�A��x.��D`(0�_��A�0����EV���i����p����'�<G����gM1ֲzx��@�0�p�c�ޡ�\���E���g��du1!���L�j��������.�E����//�y3@�̈4)ӥ�l��4��y��b�J�w�^�YJ�X�5�{���t�횐ߴ-��c����.$H�}n��#��&�1��q�������Rn]���4_��/������?;��;��8��r	Q������b������`�]{r���3��﷼�����ɤmǪK�c˄���M�Y�F��zdB������.�@:�P�ڦsӷ��6���K�BZ��+KqZL�|��~@C�Q���e�ɻ�+�.��Rl��N� �;��3-�ğ$��6��yNv(�$/t�C��}�r�6`9]�&Y�R	;4۔��Ұ\"��M����.�
�42�'�ŧ�V�TD�V��A�r���0$<.��q��C��¥Q�L����S���l�=�R�ze���OnH�s���婿���N-����ȉ����t�Y �W��Fыx|��ۼ�"+W^r��?C�G��}ֹ�E�>w$�I���H�-@-:N	�q@�a���m�ǀL��ԕ*���}n�U����(�7T��
OfhX�6�o�3�4>��$�(/-�d�ꀝ�y��϶�jݒ=�Uv:�m�E����2��N��O[zkE�7�M�&���|��!g#�*�9s%X� Tl�STVY;R`����4K���g�����4�R�?`��଎$�ɾ?=Q�Co��o`�z/J�T)|�7U>���(s�q=�N��^�p�lWHWroF'�p�lh�o��"�Ap�e�r�vb�3=b�\|��$2G>�R�{A�c�$n�@+��UM�I\j�o��u�+�O�|˦l��~~ns����`M�'�AS���� '�N���N���%ءE��BÇWїݢ�]A�i��f�|G��&���@��A�~������#��';HE`�Yd(L��0���J�*��%}�q(�m���Z4��-G����D�Y����B�����N���(�\c�b�'�%�"��S��S�0���Y�ǚR�Z���|�b{}�3S
�/;2�o�M�Jō�Kը�S���51�8(�)�F���KM��5jУ�Y����h�.�;� ��G�B�P��3��A㩓K����r��x���M-�m_b��אJ�!�/Lޑ���0<���𶸺F�AC�Rm�KY�R_p%����q~Hdŀ+5��Q:�9����D+z��F�M2oaY�X�F(��z��@t������W��߅W��<�02�`ĕ�
��[SM�>9���¥��P��\�hPIۉKE㮬����<�dȫ1�P��oc��O#+ۋ����\�đF6�PtL����~�^�5�����
2���?�iq�^�i�����9�	j�J4k���3M�iC����Y��i����9*�3?6�Ax�r���'x~$��~QG�TV�<p����Q>j�����?�Ӭ3-�ot*����'�y�5#�ax�1��8���L%��D�YA��t};s�j}Jz��.��5�@��Bh��=CƼg#�Ŏ�E��:}�Z��݁� n���z�f �@j/����hK/<88-|��]�,7�w��+����}[�����Q����܆��<}cx�O3^�����ףn#4�P֬E���{/Dߡ�07$}p�f����{�g泥]�h΂i�Z��@��ެB��%]n|r��'hS"vl@��c;W�9��~`�A�A�SlDd��SD�5?�4,ȵ�9ښՃn�'9��%FPqމ���O: )���±#Vw�d�����%Rw_@�7��=�|����W�+�PĞ߷$<��,���
a��9�ߵ���*���Z����S-�	
�����, �@���?��i�>����闌F?��dH)ò�4���s�֩�@��%~�n�'ɑ�z!%�|:X��M��|�v��`KPޓr������D�1i���Ayǲ�W�7��q}�m�������5�-P�n�l~�����"N
���c����M�J��gh���GTQ��c�'آxڌE �3�" d�S�O��ڀ��S���	H'�eC8��Q��j>ޕ�,��G���C�l�"m�hY��-��OaLX~����94�}�gd���W3���q8B3b�'d��'��R��>��\��@�~��v���ф�P�z��[��>3��o�w<��.�ݨ���<��t]�rٯi�����/	�8���h�5f���d�����"��o���AI�3�:���a��%���cכ���֛�x��Ү.M��g��9���p�O�m֣\p5ᘫo��N���Nl͕<Q�	����6��p��0[�)DWGdOja��s�Ti�e�̤Wp���1;)��.�m�0��[a�o�u
��"����38�~6K�.{��t%�`X��*uS�6"��������q������f3Z��Cx���hC���N���Vt�B�=B���-?�vj�oOHU�E<�w���g���c�����C�-fjYc�s}�?cױ~�j���]���%	�>��܍�A�ɱ߃���4O������;ɑ/��?�Н���wN�3%�[��qi��)F6�QÝ�VX��m�DP� ��@ K����Q���cr�c��&-�G~�i�n�����¡�U7[��/����^��\�eS���&XCX5���1���O͛�T_#������L�'R��д���Ȟ������.S�#�P�:�D�銃�̒�X�dێ ���j{7��~ԟ|3�?�ћ��0d(k��_� �ۺ�<"ىײ0"2#V�=9�%�g!Y[}�V�������s"~�*ȏq�hXᨋ��_pW�¾JZ�Cq���'+8
I'�!f��b�Vf!���DV��\f�(�#{�����t�`kw"�Q�'��Q��:�ho#�Z5d�p���v �$���#Z����R�0�2Ô/}�l߆�����wK∫d�Vh �PR����ߗ'_�?d�k]d��P8��L�$��)i�>�}:��0x��O<�X�~M�^��P��24 �7�o���\p%J�	��Q�^=p^;��7�������zFp@Q<b)+���Q�.�����6f3�*c}��އ�N!�y��I�� _����Mي�lW�۫��˫��`9u,�馫��?�:���O@)!8cU0��u�sW��(X�y�m�7o4�g��YA�[1�\�dV�/?3(7�G.K]��Hyխ<_�2b���d<2��N� �B^���52YSB�\�oi ؝r�PO��z�-����� �!zZ�
��x�J�]fT�(���Q�i����w��ֺ�����E�bZ<H@h��< a��[�!\ttKGZMՒl��nC�,��	ָq���E��.�Y\��6�\��~���3���W����H��9k�Ql�����S+�#�[�/�ݖt�͌�Π(�NE:�P����P��S�_���~u�O��}�[O�c�.|�9D�T��k�߅����Y�����h~���Vqh.�Qm��Q<�!1��]ק[��Vn��1x �j�f4_���}��T����;�[�����y
۸�,G��tri��l�(��v@Ԧ}v����͖
��5u�&A���z�>p��
��[���4��T��E�:2I�M���1���sA��v�!��\,瓰��___׊7�.�n��b���J�}F|	����F����2��Q�v��L���x����AF���u�*YdY�:6�L
軳�$�uqhC|}1\(^U~��	^;���!o������V�����T�u�\Ur"��$GR�]�`��(�c���;P>�8�UӮ�+��@L�o��Hu�fI���R��=�|U)�ᴷ$OAy�B��m��cvH*��w�%or���00R�j8��S�Eg�{]�aMd�F|����z^�t�\/?\��SSp��q�|ZXC�
8��!�S�z�ɸ]�Q?\ ڎ)&!O�ߔ�h#@	��k�y4�Q~e�wP���j�-c(��Ŝ�ݲ~-O\��T=�̴ʤ/�D/o�D�@L��Q�oP�L�T��)�k���<nIox��� P�Zw�l
�ӂ�dɘ��LS���(�bL.�O+|+uJ�tJ��	�b�I�
�H{��R)��i�&D�C��}��Y<@���Z��ܖn�Dz��3�18�q�_�gjQ�Pb�0�Y͞��Ζ6xWO�O3�H�*w��ΨY��<�R�ٟ;5���u�����}��H���1d3���D,����?��+�x[H��D�o��{)�~ Tʵ��i�ʗ�����[��a��O��|�Q��s�5=�\�M+�s"a��E4�V�����R}����	<Z���w�g�_v_ӻ�۪,������.��ͦ���B���
P� ���<S3b���ؙ:������n�IO������4?/ˡ�b�~��͸ִ#�LP�N ��i%b�Dӛ������M(zݥ���)�p��0Qߗ G=��PWs�����_9�$ͻ)nK^Av�5N?p�u��Q|��iy���C��D�dc��$��JD��P�!��ɼ������0�eo���j��O��*��VM���x^,�ɚ�^�`^�:3 �3��@���~l�l�%���$w����䁨2S뎓VN�|�P=�i`˃�>�/�z�O�	�����D�6*lQ���M���[�V��:�p�>p����+`;�;t���m�H���ґ^���8��i3���>��S*�sD���!��(�}��m�On��V
,$����lI!(R]��"�w*yΏy��K7|�sF5~�����<�ϒ�-aPq�����* �B9n�R��Q]�0O�D����^�c9F
�s�����ʫ�DĈ��2ʡt�XG��l��K]�?�ĮRK���/�W����7s��b \G�Z��D���=L7����Oؑ��E-�MnR� �0�V�X_�Fo�ij��Ŵ����\M�r,p� l����k��wC2M��-�[,�!���D������ߥĔE��i�.	G8ў.�Ë{X���BJ���@Z�����ߑn9�=��L1yr�<���
M�75�g5�B����R�d,B����n�?qM��!�q��y�Հ��*9�'��s��Kv��|P��`35��z$����*��N���������7��x�I*~�&S�ɜ��+�}]�ܐ����K�V�����6��e3]�K���w	6S��f�²��m��Z�T�1��u�C�KKh�j�Ԋ
�� �Z�KK�Wx��yNe"[�P��`�ڴ�P~�-O�{X����9�V�v�7;=D�`O�K��	�ƺ�E��o��[-�aY�q����^��:k��W�^�&�'+�����ܟ�I2�w$\�ޢ�����E�SJ�(����0��<�.���y��&���/����rW7������t-�.�m���c�i��"���9tT���#����N�	-�䌓+��hW*���]=��`>����Х�[�K�0Iu�8c�hۆe����1��.�x0�Il�!�|��j˙�6#��p����|"Ȅ��֚K�����
ɵ��C�"���,9Ǚr�T4m�P�b����>��@{e����@����c=�D�cRe_�ޗ$�T섊�%��En� L���j
�7񞥲�W�/�IGS���<�?`��l���"p+��igVIe"���,�!�7�:Iaǲ2��B���A(����޸s�#q�e5�ˎ�|;���r��-0��[�{P`Hy�{i6������_"���ե��n�fq��hԓ�I;�	��314A��gQ��R���r��W�}�<��T/�+�S���DG����ۍ+�p�?Xd���*�SA-�:�Z.� ������	_
Ր�-ps3�a�Ri�&pR�Շ���Eʟ�E����ۣN���8��r�w�ym��A�a;Ա"v�B�PZ� �T2��6OֶD�{�F�
X��(��  
;Ǘ B�>Ob�δ<x����va�2��4s����Џu�J_r�O\�����J\�0s��݁����6�鲔r���KD'�Y�s��cN�F�X���b���s�y�B%$�����^�j�[��4F���OX¨p�o��1��g�R99M�K�@��v��L?�Ĭ��t؜�߼b�L�(���$&.��gXH�Ъ�d��յ�ɏ�]l��d��S�~�먩$�V�$����-�����j� P��^�0<ͮ�B�	!Y�=G�υ��|I�m���5�L7��:la߇�TE���ճ�����H�o��P�M����n~gؚ�E5����U�^i��8��.8�l��}ȤOUyC��Xɀy���;��{y�Y7��p��M;V�_/�RL�B��l�#�_��I��b��F���P����bیM�}���\�!suQ|�/�CK�F��q��S�o'�ݝ0�P"ݠ�GKx>JR8������P���D�d��)�?lt�о��1��4]E�ι^S��&0��y�~��"Ӽ�~%�p���Rg�	m�`J���=��.mxM�3v��cAlb��J��w��RF�J�>���C�K�i�-Fu'���n�akT*�͢�o��a��
�>.�	��k弈�6ft��I&��p��#�;�8fߍ�������5-��W���Ͷ x�!ݯZ���J_�~Յ�k�"�+�:V���I6���@��EQ�9¾7~B����u2�,|�e�F΂��
l�*W���iu� �v�Jr��"7�v�?]�=�:t���N&r��X�6nw!�Jek�<�A��桨����U5�~�T��j�S��l4���}s�Ô�V���(�}���[Q��������<�j��5Ә^�Zx�qb��G� ��&c�Yx��]�q�����W��Afe�t"G�3�ϔ:�Y�&�Wyf�	z�n	`
Gt�������6�W*�������%�d6׾�V	Җ�������ǩ���ak�W��� ����{���Ǆ����M]P�w/EL+��U������x�(u����n1��]�	.|��6OY�AQ���b��1�ÚD@.�!�s�sj_�}��%��$�}�/7�9��jLT�
�Ͼ�T����]J[z����Q��h�}ů��"�$!�n�o���=.bKKn�_�Mf��G��$T���tiن�,+���2����p5N�@���.Cv��D*�L�zӧ�,*5��~Ć�ԃ�
۽�zn�_�x�8%�7	��P��GI`�y�.}a�×i�
�[�zά�����X�L��`���9H Tn?����%
����{��S���ߤ�< �@���X��3F#��z�~�ڏ({���BQ%i첹��V~�kq���#�K�/�Y����g�����c���������6RR�O]i�h�_AQ��?��0�!ن
�����߳�;d�7���s�ẘEN�nDyv�P��).���o�2M\$x��,�����!�v�h��Q�Pn��0t	�,	*Ɓ&2 ����l���Dw2����S�j9e��/�E�-u�/K1l���и�S<X����-��I�H�����/���.M�� k��� �J�HwUҶ���(Xb�q0�	l�x鑹���Kתq~h�� )�'�g�B ��lE������fR�h�m0��������C�G�M�f���<K�&����7���J`3�[���[�����A��m��bv��1SU1��U�VM��K۰Bç�hҭ��k�N�tO�.�ϼw���?�t��b��4�N	h[���^B��-�'��>��@�g{��v4��A��{ KY�(H��Y
n�#S1���ԫ�ۆ8M<�̬WF�����
!����u�\h�6�X�7��@�I"˴uW3�`��_c��*ˑ��1ߟ+܋Y�*y�����.�y�w6{�ڦ���S�"4>�����?%e�w�K8��=r鱍��p�a�����ą�(�<�A?��eH�[��msL���-|��q�OL'���3�����T&�@���EcVϟ����:�Mo�Hw�gށ�`R�T%������I��ե�%,�o"�]>waP�7�x��~�,֞��|����|��J��G�����e��s���{������Нj�E匣G��'��8o��2���^���M!f�n�v&�}/z�\�DZ�LG0hZMD�C���P<�������Z!��e7t��ه����!��	N�
��#e���,�kQf� 2��p��穎t�A�1�*��3��|}�M��Q���t�xx汇�~<r]�׌���("3�d�6�d�
;�4 ��%z��{bȶ�-�,"&EÄ�M�1a:�!����gy���γ�v�d��ܒw$s,F(���9pe� �Bϒ�����`i��fz�X��������醧����:�薟�������f�j�[y�����n�]z&�JAjc%Ј �Zo�/#x��/D�@���oTϜ�5H�Χ �`�ŧ�	�VL��vF7Cz2�xyL�G�ثY�̅͑-0t\v*����s�[�t�����h�i�^�]�7���\y�����&Z�W��{�c
����qMS;@~�m��%N�	���h��)��uѳej/�M1	��t	KnĪ"��W�^���$����͉�qަܨ��qZ�G�r��im�Bb�V�\�����>��m��U6����j� 9���r�8�$��CF`�^e{���S}�k]�/�G���'�I��s��Wf��i���jU�P=[��S��߆{�Q$�ݠ'd��t��)䰽S��w-��Ð����Y`����_|�C`U�8n3hLS��!Pr���g���}C~A������>��[s����-&JJ���X>���g��\:8�R�I��CDW��c��}��}E���F%���HI(�>ȡ�P��梅+0?��6��Ҋ�]P⥾k$S�a��F��آҖ��h�sp������llڛy�z�`���DoP8�z�f$=��`Ey6o���~7A]�R_i�\�W"��@�j��$�qpu $vj����i�
C�԰!��&H��<q�ꕈPf��@s}KփB,�Q��͑�� 1�c��Pv�%�1ʅ{��P��\��6��]�͏����T ��*o?V����ť��(�񄀯a��	��ս�H7�T��4e~G�ӻ8E��M͋@�Y�8�(k�Q��,���vM����~�'�)<>w��5��焄( B'(��[cI����B�z�Z#�����}V��a�ޖ�����|a3��j�2G��좆�.j�vl^�Lz�+_�i,��NM��Y�!�Y�V��̾��4!�S&���fp�B�Cy�S�)C7k��� ���j�!vt']4a�"X��/�[���m �+e� �ѯ�[8&	
BZ�4x�bϗ�	�߰<�s��ʮ=�g2�������Sꇊω��}�b�)��Gg���kc�TDq�=噮�0.$p�����H$	��&Y>F�6"��Y�4���y���e%��.LԳUm��X
}���~���%s�q�3uhaȹ��ft��]���ރic����T��">n+ܿ��Q�z�5s� �`Q�V����%�=��wt)?m���;�{�Yl��MP(�P�͖������5 �z�ۮw�gDfߏ�F��T^�7r�qzz�����R�L����kn��A
��������]Q�/�e�-9�1���\\A8k�돚 ?��iП`T�����(I̠���f�zK���.�Dc���J�2�[2�j����h�#(�k�^�%�Ԥm`Y;I%�@6��K���ah��Ux�H�Ym�q�H�,]������理�m|�e!�j�]]r Z
6�)�����rk�кJ
�x���KDȴS0����-;����n� �Vl.�(�J�����6�-^��ʤ�}��taB����1)�o�/ԡ�E����(���~���P>�]Zh �=��Gh�"b)��&7v���@}k�fs(�Ʋx\���J�B��r��F�ܵjHp�qA��Χn�C\����?�0�?v���i����O:B���%� �XR�I�^C:��g(^�At�03�z����u�u�{%+�m���F������MU��R�S�])n�s�ʮN���'�Ȋ]�o�@�K1���.,�n��\����Xuر�9e���G�{a b8����[���)����VU���&��}� ع�P��کk����h>:k�I̃f��A~�$X���*��#D�r�@� ��2®�'�#�,���L�ېs�BY�z6\�.��\�^sÃ��e����,�Z2�9��
*��P��xVM��v4�#�)�s�i+Μ��\��{�m�ꢇ��q]�.�`r�`��"�h��%
Ԣ^�#���������B����W��Y�-����^$N�_p�qm\�n H�O������HY:1H���v��1���og"dgu!����@Ԃw�B21�v��f�L�Zd !�E�l���/D���Ŝ�,8��Y�#jϽI&O8*�)4Nu��$�ؓrUh��p������k��h%�)7Rf���dXS�m����"���x:��uERK�[g-�z8=�)������/�o�Lab�_�q���=�t'R��wߖ��_u����H,u�E������W|�<9R4��3f��R�\g��T>��YX�����ƋAǛ(���O�t-~��'�s�v:�œ���蔐ɽ�.!�o���O��S�$�\h���.'��P��:��,�8��a"A�nT7g��||��N��ip�u����O���N��DK�A*HQ:�T
���^n�ȶI}ͥtY�0Q�/�u��Ta�q<Ԥ_6��X�d�*�%�BY�h(�ͯ��U�2�:o<��y���cݔ���9h� �"�r����)�p�&:DKϾ�"9	����i���V��PKC%_aq��62�=���	!�9�>��z�c�*Jݭ�6ETZ���_/���~}(/N�K�V�͎����4U���"�ǖ�"s��Q�0<����#���!�2�ы�Fz6�U8��;k`Z�	
�A)�c,�4���jG#���.�U;Jț$F��<��,�=�'W	�F�>r���{�^/^��~ Pqe��$����_�6V.���g�Ȇ&�Ur)ߞ���ƶ�>��(_��e�����W�@88b���2�s�P�)�͓��@˺�N��*�~x�o��;|B���II9����}A��0:����^�/�
����,�/��3�>�h�M���?ƌ��ł�V{d�qW�r��UZ)��}�+����P��ӣ!�w㰚!%dy{����t��"��`U7vś��9>�9h/����.����d��&�l����ZF�X��2'�|0�I�/lLF�~��_�q�b�9��}�q���J	f���<2��2s��y]KbX�f#�Ƈ'�>ɬ-��E�NuCa`�B�A�}l���#�@�,Q�A��Z$k6W��?X��T0����_TM>�~2wyn-J��Ěd>��7��u�g~��j���2�U.w�x�=l���<mp�K�*�4y_o�'�:�a3�A�)���&�:�M�+8�Ie+(Ab�)!�����nD�)\a��9��NFk����D`���&-�H��S��|ڟ�߿y΋�5��d�Sb\-h&����G�g�X=�3�J#z0Q�N�9��]���m�0�4H�Ì����G���O��:��
-����^���O0���i��y#���壣���*^�h7���d+_/dCP�Y�=��-�(��������+��{o�ݢ�n��rf�#9\sU��#.�B'~�V)Av�xa�"x�ī�_a�Ⱥ���X*�2l
��d��\��O�c��L~��U���'՛1fC}��^�T��#����A��H��G%�2�YMFjG��)>�)���ƣ�uV��[��沭ۚ)}^)�)���t�%X+�a��e~�� ƶu�TKI108?�b���'�U+��j��@7� ;��#�V�RK.�M�ZmI�����hJL�ʈ� ���e2����(T�J�B�q)v����l�=4~��c���L?�l�H	�c�����$��z�z�8���7�G.���&�M���J^�	�CF����@7��B�����^�`&3@�h� O�_ڼX�:���3�W۠�RSt���*s$���i�e{�U�D9�b�	�S��Cq�rXդ����Q
%mK-�˭�A��E�������BOE7�� 8���) ���]�Il5֖���X���{o'��uCq��_�I�]7��f���͸�r�� IA��ÊC�}&4��8���j(ы>���"�u�DwE�|mf���V
�²��R�h��֣E�+o�pw�j�#�DLn�?D.���f�	U��f�+�jw���F���X�I�QRݖG��E����-P>��$�[$�z)�Ɖ���bN�M$��VW�o&%�C��g0�j�����"2���V�N��gjW���������]���GD�&_�=?�����z(A~����%{�Zf���L�����T���eAao~e���{V��Y�<~pHm�����<8q7$�.���\V08�^a�7Q�wZ��q8�1�|��\��c�̶���8�O�>����6��9�V�'b����)��p�N����_#���e{��)�����Q*,��9<w|:9*��[%_�5V<�H��Vʢ��J���w_��5�$Q�~�}%n�D�Q�Y��(�݇b��� �K4
V ;xdl�{t�ûk�}$D;��c�NL���!>'���xR��`{�,7+{C�sC+�K��q������k���D��4�+�W%8j�4u�Z¨q�*��n苷G/cʝ$�;t&���؇|�td���|X9�z(	�ͭl�a��0��m�Y�� "Nc��<m�>�&���B�x��q}���/�?�� ����uͱ���p#�ì�tث,�[�Zm�2{2��������R�N�N"[el�0�%ck�,�E��WS$r��-�@�M+�ʴ���B�X�A��P��V6�8^b�
��c�u�"�SHXk6͂����s^��S�xIUh'1�3AXX�$.�f&��X�ߤ.��P�־C�
������v��V�g��7ϝh���#���Cx%��4>
Tg}&�SH��71��嚐Oz�(p`���Q4���'~�1��2.��I�oz�pl����
J/;���t6ӣ��k=���C#p5O��j��[�֭wD����>�`�T���]���c>-z�6��;[�V��T7\:h��t�"'����ظ\�h�1�u8ढl�B�u�����22���A�W�n?�e�^E{�YkE�}8�J�R���z�]����13�����4&��mH���
��\c�%�i}�Ե����j���(E�)=[r��)�f�
Xi����*d�}p�g�Um����d���a�(A��#e�O>kX��/�ڐ+��̙��޽y��z���JXd�ϪEߘ��3`mv�K��|7ʹ� t�Q�	�o�'��QE,��0Y�ɔ���!t������)߁���(Ҡ��=Z|����t+�6J��dE�-��7`Ť!���c���Nh�p�|������̇�f�����"��i�����:��b�'ˇvS��Tu�m����O������xe�)�W���V1�˲�K1���z[^��Qa�^K[v���Y�z@��g�1�0��M[�P��n��9�K�Ϟ�W���1њ7F�O��X���S-@'��}Z��5χU�{e!��޼�O�|2�%����H&0!�Wa�=l�2a;���`���+V����yvs`�z�=m暯�Xm?���:"���4���\:�w�/���[͹��F�;�'��AkȆ��3J�qP3sh������*��	ͳnkQ�E4F��"��J��?�q':e�2���U~z0�s�օ5�,� �w�������3�����ED�������&����W����dNX*F���-y%<�l4���pd���~w7�4��}� ��sw#�P)lG6C����c�^�X^B!C^��4���b�R$�w���o�b�<��<�Ͻ��~�G�Փgk�j !'�=�Ǆ�0��
��+��+�2aÊX��B�G��>&J�]JVE}D#k�\?�f8o�l}'��i��r�'���/��6�B��W`�D2P4c��d@ҵx���`m���m��^�:��F�xr��� ��d���.����E�KJ��L��~B>�'��^���M�߳�r�EXN>�f�^Ⱌ\�N� ~�g����>Ͻ�!���ɘ*ș832��q�~6�'m��"J��@U,sy�Zo/��q�_C��F����!����HB��W=�Q��<'~|�[j8���/����<�L����6=�zJ����i�(���R���S "E���n,P�L���2:l3�po���P-�$������z�|��C؉����'T��j(�kI���%G���ğ�8�M���#ݬl|Vgdm�4��r��Ra���M<��T�ק6�o�U�8��Zސ�o�󘖶�P��A��N~�����h�.=$x�Iq[WI��,n�I��q�R��{	�ʻ��H�b�5*3��(�5��>�>Q�� ��
�|�u8�[�b	~侸�Df�_��$� ��6_��L�Y5�r�\�`c'4�8L�2h�'P��^���|A:v�D�|$�|��\�5��S�� k���������[R�U��a.���XW�hh�Q�SG*�%��àRJ����y������?vs�ejȖ�8�F�[
�8��JHi.R�i.��c Rm�L��y��A����?;5�?Z�G�����H�B= ��򎈵�g�H�%��"q��-`�-Ǹ�]��t�r��My�( ̡\~,j�VL�0�I�hd�m/9�����V77�ۧ����D��D��E�If�]�t<�m嘉�k��D%�w�~x�>�N�2�2��~����d�9"+j����D�&@��#���V[�z�'mFcՋ�uKX@
�ڲ%6������`�3{�+��X��2H�e=P�����C��G�텡}�'j��N�>��I73�iH<�T�6�d�������>��xy��ᵬ��zTq���ԑ�����Ԝl�)�:D3x])n�������l�cv���jc#e]\�?'����uhgT~���L����+d�S��5��P�@(X�69s|�N�e�es��>����<ܸ~��e��`�8�Ljۦ��0Eh�����)��n)��1����Aj�~�M�zc�~��9ď�hJ̗���h�ME����=؞͞�z�
��B�|�u00�*��
:Ԣ�� ��L�6 ?*n`\�.vPR�N�6z�tqC	����o�����s��mO8x/�v+#bP��ph� /[g���[�n�Eiڸ�֖���G�y�
2�C[������zº�����5���u����d3#�*ɿ��k�6Q6�YZ_�xAC�br��ݣ�;��%Yݛ���8g���"[�Ifd��u�IJF�@&ŀ�M�
��Z�����Ԍ�Ϻ������a@ ^�i����rW�A�� �=j��I���z�MƜa�v��G�H%�F�.�9�,���P�t,���q��'M���%Jn4i��EwP��>�����V,�P�5E��تc�# ��g�6�߯�m��;���jP�Q՛b���i:�|I�)1�Wh4h��S�ǧ$I���2�a_q@Dv�o{`O3��d��N.��;��*���V��A����s��.�Y�J�G	�%�Y%J��WKyMXf�=� ҋ�{\��[�\�Df]�_��k�� ���Y���$�g^�x� g��i��!�#��v:��Ss�yN�m�|y�6>�+X?�A]>�I��S#$ө�:�f:a��V6v����zc����?Qe� ������ZS��z�fp��lEݱݞ��G��/�sF��B\Cw��t�Ѥ�:��
g3`Х"�ͣG@��E�Y��PA���G#P�8��/�r�5i���}�w���{49a9Ay�y�,ɅK(���(6)��*	ȵ4h��$(1�05�ɿ� ��̈́k�>h3�FfJ���^$�u���Dl�j@��g0@��od�/��j�fX��CAy��c0�]��qĺxd�����}
��?�1ۏQ��h�Xܕ�Z�#O�e�&N�)5�,��	{2�����J�C&1'_�A���K[���̀�T?d�?���B�^���5�ޭ��u�T1�E���О�*������������%�i9��0�Irp�Õ���I��bC��D�luP���96��l�;@p�w`����|r�N�r���\7`���5��}�<�z��x=8�̈R`Os8:����<���Xh\�#��/m��w�69sn�>�L]4�����o%��
o���jt���_!�� g�z����l뽼w�	י�g�E��G�D,�,�����Pw�k���]d����k<�R8S�w#�`h0�DH���&�'��V.:���@���ie���{�X\���n��\L�IJ>���d̻K�%�G�q>����u�=#�Z� r�ZW ������e�"}ؘ���&q�L!ߍ���Oj�����ֽ�W��%?�{^�|yO�!9���u��/�s�.�u
�8G�1�##Z��7��	�E7��:j�'�^W?��S2�h����Z
��oh;�g�V���x����b��g��{n[*tO\�Q�pa��h�6o��d��1�$��n��)&�� 2�QqEf�ح"��x�\��o��P;<_�q�l<�(��R�����B΋����l���i�,���v������&��ʴ��� ���^GGbm*�h�aV�8������dQf�$�p"ޖUv%�  vC�y�qw��,��'�J�N�k���1~�Ψ~m�ozAߏץRݒ��em�3���^r;/���h��v�����M�;�W`�B�3,}�!^��@��vH>�G������ �¼5�!�C�oJ������\;�۶��Ä�"�Ş��11L8�W7�Z40#�/�L���pG���>kX�7�����e�W����v ����Q��#N�6G��J�t���y�WřH'E��zC&_t�����s��#8/Z3�*��3�@��Ԩ��#YmSK@�a����wB�P���0j��8�~�ub��U�G]4I���M�X{F���46e8�ٟ�&*�Ba�u L��2�z�8�<��(V)A�+<lH�	�����q���?�����)�Q�i��b��>o�Nێ]���E���#ڒ��}G������J�.4(e���p)�釵���l��$��9|�vC#&"q���K�!N,���B��\(�й�"������fz^�Z�)ݘT@ٟ��9}7�ʜ7���	��$���6xC�nT�=���!�q����.m��j���o�i����',���j��	?�������/DZDsxBn�%0����0��v��@�B���)W��hHK#�qG��/޶O���w�VL����y�q	4�8˙�J�j�[�+T��C�P��
[�޼J�S8)Tsφ��ך�}2�$tGn�Z�R�dO�} �{�+���c�-KхV���ɓ���L�\<��_��׎Ĝ����
 �<�ȉ����ɡ@T��Ə+��_xXYm:��%ύ�7��4A�D��ܲxWt:�%��sy����dI��b�KG��W�'XPi>�~��
�&˙ ��\XaBUO^��9�,C�B��-G���̆����f��x�ϗ4��ā�F�'#4���Q�_�#�|@�5ȆU?s?��Nq����?A��d#A}PI��Uk"&5֙o�զu{��5NIp��J��������>\&�W��l2;L�Y*���CG1qSb���*�X�/�u�ge�DO�B�F��:I9Pܐ2Rt�<g{~�������?Dl����l�[ ޣ�.�u���ǡ��~�ތ�hh�(ꜱg�\���Jg�r�	4�ߐ�*����N��i��MgEIHU^�������'Q��t�qqү���]X��{κ�ԥc��2 _^T_+��@�z�C'�3�!x�i��VD�y��#9�1?���q�s�*ύ������)N��!���B G���7\�FK�B�!Ƴ͆�E�������6܀�+r9:�:���%�Ԋu@���4[,o��,�=L���>=8�[uʪ.?���$�,%H��u)]�ٔ=n���Q,���-jĻ��14� W��!�_���]kg*�z],�n�z�W���\̜b�BF��$;�7�|��|]���߲?%KrQ��hu�2{��?�4��*ʕ�ޯu�M��9ݓ�
0-jZ�5�t�q=Θě��0�-gV_{!����y��i�X���&�������Q��H-}��DR������J���5�q�߭1�R �qb�;��o��&ɴm��w���ыp���jƖG!<�K˝{���侔�D.��t�����Q�q��^
�4 {݀�:E�����9�夅�N�X�X��AQ��ؼC���Qlih�'$ q���y#�7"�Hq�Y=��k��Bx��e&�|��g���T}Ny�Q�)�W#mj��ꧮls�����U�Sg�x��η)�l�R���댗>��6�c&�P����@Z���ϖ���VR?smP[�Tɥm�:�z���Wy |�F��}�����=�����K���J�cAd�i=��ɏz,�TJ+��%�*��R���1Ƌ���s�6����@��>td)�����+*�FU������B��s�ϭG����'蛧G�53w�/�R@۱M�I���i�J�c�A���\F�7/36�"�w{]�!�}�'���+��X��@�Pv�ȿ�F�D̖��<ڹ����0�nM��]�j��f��3c�CR)�'۔);�-�
l6w4�t��H���y䐯��?2iIᝮ�v��#��o�܋�$n�!�\ÙB�:�����D�ߡt�3�"qi|Wwkм�e��sW��O��wҗ�1U�e��8;�$�|��û���ګO����	5��V��xuRv�0����X� �I��M�f�룈bT�	�>}��-��]Y�X��cp�������5i�R)]Մ@���R�ӫ	T���^ks�Bp����U�.6cs��8�Ǹ�bqO�Ro��!�Y�r�~^������3޸$��qn���,
��#R���ѫT�M�ǽ{5xj5�?6-Z	�>�Œ��N�|b����$��do���c�Q��E�*�ǲ��b�|q{��}���������Д!��E�
z�a9��X��W�۰�U�`�r��o&�++�Ol�=SmDQ�E�ѵ���Z���ˑ��2�"Jم^20�LU,O��#R|jf�g�p ��� ��ga���
��e���s��F�E��|��8�W�xt���'=���j>W����х�v���g�O�M��
��*.0u92?N�"��L�RWKN<��B�> �]����9����.���Ԁ�j��}� t0�H�֍O�NUck���������u�59N�`<������iŤl��q����=X%����Z!\�_�0Vnyc�)���t����~E�\b�S�� ��dHX}�����c{ QD��\����ںr􌂲��F��k�~���(�Af��ؙ##}'��JP Gs��\�:��@���n�#�Z��y8)�z��E�MY���n�g�K�#�GMsr���L?l�f�Q@/F��r��sEz���1����Vg��:x�u������2�5b:�t��^߰If� |eZ��>s�����+BNET�(];��Ì���}N�A��c=E��5� �j�^eD��{'��e�xchƬ% ,.��;�g�ӷP�QK"��) ��n�o���r��\����ݮ�{t�f�V-";��2�V����G��������Y���`%���rq*�V^�ճ�����g����10Y���_��-��3K��V��=�ʔ4��6�\ԣy)Ѽ�x�]�������V[�'�(pq�	��0_����x��Q�P��7ZfwU]���_1B3h�T�X��t�L��=��3�z��V�I:����+WKZ{�ho�	�:�=@P�`�S�Z|uK&���"�rG?�q���R�E�{Xjh1�P?�B��/����v�b��XA�bQ��5G��P�t���N�|�˙:�w��(��
��TL���5����rf�s���j̎����X�a�clؤ�%�A��jp�I���>.�Q���&��8��Du]�9���|l���	~n2�c��Yա�,a��LR��K_�r!;�Z�'38��:��Ф���x�a�ߑ���!W�7�|��;Dے>���:X(�Y�����j�GY��h��{���qs����r���Şr��A-��O���0�Mn`�I��]�����K��r���~����u�$8�xN�l����S3�Ek}��Tr�o�~��̸��ڪIW�����!��܉����˪w��"0c�}�V���hD�N�Z3��fk,�=�;��6��U2$�b�4k��}�T�,�`���g�R/�p5��mSY���t� -5$�T,ρ����̥�As���71s)
�^�[m�@d�F�n��7�P��[�F��^�wćد}Tb�Y�^���/ͪ$�|9)cb�)�t9v�,���2&�포�KT�,�"@�L���$�\�(9�GU�s4��2e^&"�y
S
���bks�~J���h�1/d`}q Sҟ{�Ҏ]bXϱd�a������l�=4�o�U�T���^5)6�\(tq�B�8�L�4֬�J �_��=�j���2J��>m�̔\�Mb�Q9 �)z�8�
_~����g�|_�.%���|�����2�C��7�,4Z�����.Iذ��V�h�d��c$c�]��Z���no�0�-�B�i����umL#��(8_�I��l/�y4�U4w�
�I�@K��&�+�ۻt�1J&6����Hd�) ����R\!��5ix�I�[���Ϙ�l�IXH�y���O���ɂ�s��}7>�'�w/�6~ᒞ�Ҳ�5
�d=�XK@n�g�AT��K�"b���%��%����\t���p~�=#�Ff.s	N̈́R6�$F�ڲ������ 8�y���� .D~�岡9sRc�(�&dW��I����T�3(^��Ă���ueψD�8)�v���ř����(:&x�kc���X2��|RfM������"���Ȳ��Y"}U���+����R��}�4��-__��Uy^z	+X?�^Iu+�Ō������Ŗ�U�V߮��s�f���|�B�	�ɑ������1-?~�b~���ߏ�}�(�zP�=��e�4�)o�Q�'�LL�zޅ�����O�3H�Y�u٣�۫�uO��Oܹ
��r�+I'Ճ�'` ^v y������-�᫆�(�0���Y���f�d��0�T�ZbmH
�5�l�^��`}��!+�?�q�X�f����&RE⊾ǳ6��Adp�eP���~�"�w��w��~0u�h,�H�j����R�>S�L�D��
%�\�h������b
A����ىb�&���SIٝMob��d��
ڕ*��d�gk�"����"v��T�A���>q�C3TJED�ӏ~͹L�v��b@(_Yј�7&��h��P1W�j���[�S	��`E]lKu
�N���Rl�n�ˮ�T	�ߪ��c�b (��r~0�Ҷ�hNU���?��1�uyFi5��:"_�bKT���2��'����5WUh���܊�n-�o��YR��q����^�TZң�1�Ѽ81ޓ�{!]տ\���hA�k�F^��	g�-��o����YHț�߄/���8t���w/�\$�;e��=k=���| )�v��4q���y��,�6Z�9�G�\��������(�[2��|���`�tEθY� 
.��ἑ�+!�ˢ��"�Mͽڼ�@6��s���~Z�r7|���񶝺n;r</ ;yJU�o)��#!i��p]�[A�i��$�Nð�����CJ�_�$�7�0��iO����v�����:��8���:y��Ľ���&�A�#͑�4�5�j%�g�?��ER�.�5��,��(V�ج���7�Re�d�A9̍5�z�p���Tt�(�u�T��Ν�?"8�zm��(կZj�amQ�rW�w����m1=áb����0,"6���	n'J�=�1'��\+�a�S1��Wlm�\�IG�h8�d冋B(_��zED���1c��s#��90�x���;[Mc�Lw��[��_�ۭ��l8�q�;��s���y���p1��i�����.�Qv�v�jأ�L�a��;}���C��LФJ��Vl�s������:�mi�,��H�7���#��6��4���1@l�,��o4Q�Pд�)�zbZ�൛d'���9j�uW��~�9l�aU%�k��3�]
R��؍��^إ�Q�6��{��.2��fx-��I���0������������+��0�	��寪��?�@��l�T@P]zCCs-��e��^�4��O��$;�۪|�c�Rq�+5�}�C���}e�
�a
i��Nči��sx��I������nM.�T�s��LSv᭧�Gk��:x�Z�$�R�6h�A��~�����0J��������������~*e���Y���K���J�r�&�֯�h|C�n�NU�Z %z F����v��Y�8�~��:^Œ �/�9�ZL!}M� )կ_$$���@���U��wI)��DQ9��;�cFq�7����qKښ��T���Cx��\�l��u���FH�[�]��F:�x��U9'ݻ߳K	�L�/�N;�l�W��,ΰ�Mȳ�)@F�u�ڃY��B�K�r��hf�KM&!�������8P� L�$-/�t��J'"h�.�K7�t�k9U�Aذl@�_ )�fpQ scѮ��Ͷ	7��w��hC�j�Kl�+f�8>>�vg/�w��@�s%7��]_!v��Z"$A�)��>�}�v�a��&� ��#�_�Ar�9 Kv�Q�Y�ơ~U��]�]'�_ެl@.X4��kihh��Ve���/#�}ER2�[b��<����hcpW?'�sj}k��ht�anmi��E[��?�$�(�^l�th��O '+nᾣ�������.g,r����6�P`�n��\5�b�G��R~�۲G}���a�^y�L�\-,���W�}������bw9�︿�����1FFe��Y��NT��8�~�A-u@����QJ�[|'���O���,I9^-�>=���:	�n�]�|�˥̲x!g���=n����ɘ&(� �-����K�o�>���^쮬����D	��:C	PQ|����6�P�j��F�̌	hr:
�n��2"O����1�NKP鉵^|%�$@�Px�l@������gY�;�r����<�(_����-{��5�k9�љ�������W���H�0�eVO����	c�[���U������e��Þ��k2h����{�� ���b����b R8�2W��Y���_o��˶����F͒	�!��ő.���]V�|}���+P�D=;�|T�X�Q�ZcC�Ų:�j�(�B�����,ё�N�9��m@h�c)��P{+�ˍ�L#t��}}#�j[T[E���W����M;L�j?�P>��&4y�o��YnR���p�,V���΅��c�I�Ы��u���eT،�'�r���X���)_��}$�=Na���qy�33҇�;�o�)���K��W�i�)���}z3�[7�|�)$QWt�>Ǡ��$*� C�Mϧy�nwO���ݚ�>��a�H���pn0�u����s�U�$�y��#G���=���ѕg���,�i/��R{	V�z�8��*��Fh���N�X�F�Wb7�x�?��2�j�Y�l���������MfZ�.Iq�/ Dpq�I(V�7�nFI}�����6;����,#93UX���l���n�^���L��^�<s�!�T���?MTo05�{�&�g��n�g�c�Y�W��|@�#����)l�D�%��s�F%��gq��u��4�o���x'2M�Z�l�/B���ֈf���ȶ(�6�A�2�I�C�!���k�/��:m�W��������6��+�m��bf���@����}�g;a�K'�x��>r>Xd��v��� $$tk�i'�zG�����{
@8t8� ���;?�5~z��Ef��+Y�C(���բ,���=��Ք넬��{"UqJ��kS��Sݟ�,�w�q3ڨ�Z{� g=v;^��U�6>�>
�
�~����'�9���İ9���mw3$xb ���
T�&R������Y��W~
�\���q�ϼ�W��Qb��$�� �'\*~?ؾ}���8�E�D䔬�a�{����Q�Bk7c�[��p�<�wlG��ܳ~s\������22Z���ۛ��uj�ݸ�ls[��Hj�x>� ����殡b,.7Ъ��W�L7�K����pa �j�d�63lqU0!9����nN)�nsI#Ӈ��JFX�bi�\۱E%i�y�"5&=��f���"����$�ņ����Q1$/��D�<�v�p��$
�e�p��Ո
���� kԠ��������W������� B��w�3q��t5�8#!Ed����bq�b�\CGb��6�������?Z��3��KZ�����u}?����,(AhE?j#7�|;,�"���M
(��Mt�MG1Rp���T�����$���4�Ate��A�G_�^1��)еt�rF��;�&�7��"���CG
sy"~M���[�	P����M4�v��R|�����j:�Dn����-������[�u���͒��L��A�_�\��0��� �������=�Y�2�B�1aYb>����!䇐H�|y^�܉�Fɨ3���Mڔ��[��6�����iF+��vZ�>��1�o�6�x��g-��9�SE�F�E���[+���n��tJx5��f��y�|��L������kLP�B�^�.`F]`6f 	Ϊ�Y�]{���@��x�RN�L���t�w]������&B�P���fAU���DY7m	}��?�QbL�_o���m��~���gt�9�d{��>e4 ߆�rd�R�o=���N��k��c��c�M��tIOa�+&�M�����2���.�E����ڽ:�Y2����z���GQ�P�k_4)�=�O�C���갿� ��V���oRŏ�.:�>�t������z��ZG��:��V�s>x�
J "T�o�	W�9�/��Ɂ!�Y�����L�@���, ����D���6'T���9����%�)A���wO�ҭ:�锁���N��>,K��8��	�o����:���.93$�
-��Jï?ײ���)�65Ϣv�)��;tV�n��|,��%+: �|�ܕ�v�c�سz^�thՊ��;K���o�n ��=mCLv�D_Z��g�(�A����}��u����U�@�X�$�C���9��a�b�"���9��5m���%B����%�M����m>��e�֞)��1(v��� 3D����xӖ��%>�-�.���
fe���Ն��O?S�)��l���յ���.lC�W�Ҍ�����n��2}]�����Y�>�Ǣ͓�S��?��5��xv�O�G�*s���]�~K4OF��b�B����%�6֑���f��#h����j��2=�\����W:[�0A����@���P��F��{�Ә^���1�GȺ۫�F>��-ʀ��1��D&�h���&0���gЅ ~�юQ�'��&�P�x��BTO=�2<�?xy��Ì�cy��ȁ��3����VMt�	_�l�k�E�Y�2x�Y}R="p5��`�8�0!ˊx������/�褁%,���� x�cRãg	�����D�C%$�d� ��%���g��%�����Vbw�~��3�<W��hyf9�@s\鮷tV�( ���X�R;�mY@�J�>*J�Z��Z)I^��o0�'u"8>�S/~���1�������6��\Th~.K�]`��K˘��&0s����&�"��膇�����(�CX����-���4�=39����|X�Qҽs�VWɳ�+�6��F��t�ىq�NR�8��i�<X�ς���۔VJ�L ZO��M�˳�ĳu��@�����[c��U��Y4��w�`��7<O�h����ހ}H��ӬA�^U�/��ي���K���GxJ�&�M�0|+�A�+ ;{��p>(��MFG���k�O��^K�YB#m|�h�#��Tm:�u��"��`Dȷ2e)�WxD�9�?����J�=v�F%��,֚�񫕡����r������~�W�G6V��#B���]�O��>Nɴ8�U{�����Ҧ��w뜣����Ou��rWt)�;�h1���^C={[�gYN��ρ�� ���W�:�����B��̇=�6b��(D�hI#Գ�j��ğ`׾-��g�)YU�Y<�D��H�)(�r<(PG��V��G��4`T��^��=����^����-6�;9�����r�	N���W�]��W���W�0�1�z�o�X�Y���/\3#j�k������%-���/ J���e��D���x��3T�z;kךAf�T�Y�%hz���e%óz�|-�r7m��I�fg@��<t�A5�X�V#gY�^]���x����D��lXC _"��n`�XhY�z9f@������7:P�U'k�}Ƶ0����?�j@1��h +�����Y���&&㗽.U�uU�歑c�T�S�*���K�Gf���S޷������Q����ʜ�N)� ���Xl����1T��ѥ2��7�/sm1�K/�(P=�6I>(�_&�5|��n�����
�KeS��ً,�ylM@�,�\� ���4R��Sv�E�;" ǋvŹܜ��B�u<Ճَ�Y��^�g.��u��ʿ(�Y�k���>���~�GŜ4�0�2�>�?+�)�S�l�a6�K�R�WJ� �N�?G&aG��Û�@&̿�w�,�^�e�o�r�]��/8
��K�G��֙��<R�pC���C���i�����[�6�ʝ����:ATr��w��gm�yg�: 
����~u*G-'^��|�&�\6���v��^�ZTr�v]�9$�9F��}ۈ�ףS���+s�z�+lCm-���lT��CփF�u�BG��3C�	nt�������>�u����xԈ}`ڿT���+҉&��N�eQ4{�qq7�N��g�" -��ӄ Q��ĄPf�X%��1� &���Eb�K�g�0�H�53J�K����:��N�F?T�:�1����?�������;V�*���5�sk̂� ���Q���į!6)}~?+�.'���\����X����j>���b?�z�>�ҺqE"I�4 ?h^�tBӚ��D��'�骊�HB�u�ajb��TTۏ涯�^Q�P[o��Ry?�0�uAcoU����<F"����Q�z5�G`������kEF�t��Y��.m��Ϧg_�w��J�7�K�wkS����0�2�0��Tj!T[�)�9�b�|]�3LF�Mdt��o7S+�ɥf5�l��^>,3���T�'���� :��߲OW/��q|۱ݢ��5)���u��\=�a�Ѵ�2Cة�)���n��������E��89ӯyŭL.�{ٮ�Z����-_Z;��g��?.���o*�t�1�O \!OC`x*�o
�a����c<ؘ������ų�1#\����Ō���v���hT���������bѸ@i�FH���=��C�	ޣQ�\¤�O��]�`,����gj���a����K�c�d��֒(���
(����&�-2�~�3�x�>��x����BЃ&�"X˰�yH��5��n�5��~a��q5ƫ������Q�(�>PSed:���q/�e"����)U�.�8��{_ϐ��e��d0ð��h~����l�t!��$^���h�n��ܕ�X�
�j����.{:�.���,¼@B�Xfut��e�F�)��"�r�2a[>D������`ey�m���`���<�rܵ���'N�¦o���j��8+���x-'�o��"w̍BA�i���g��z��6XR��;���-��T9��g����/gN�2"O?o����:4xZ]�a��R�|��9�3���DD��y�v�ä=��A��N�uW%@1������)`��nw8��<�w�̩@����;ֱL�b'꤫fL՝A�$����+��q=�Cv������t��-�W�����#��]��C�Y������`��صy
�U�W�s��(�%������lY��z)�b�1�*QkW�(
i\��:>J�k�%����*�P���a�n�l�d�����qa\��2�'�URf�1YL�zP�z��p7LG]ߵUP+�hղcߦ�ca�.-�� k.�i��,D��(�{����_vwl�+�t�W�!_7ڔ�(Zď���Zi,���)�����8k��L�����c�Uc���p
��&�΍\GckGHy���O�U
:P��Y��o�1:���Q�b�]c]�+���˾�-�ޡѲ#z[W�&<!�h5�"��=�5@��B�Q��ߒ�r�*����rfL�D_jV�H��i�VQ�"(=<��;JPA���ϘA)��K�j��n�*s�`갈��^"�{[�
�:-္��vM�A&���Ҝ�HMK�ߣ�:�M��r�x�3�`́��϶%�:�ނt:����J��(���L��N�-��66V��<�V��5e����5WE��qh���
W�T���f�S"e����ޟl��)�w�jG�ܱ���G�}Q}y���CV�0S�O�	mi�=d/��"�>#�ǦХ�&��Ã/��L���� �ĭ�m���Ò��GS�gTq��>�x dI<�v|m�P�3�9��S��	�H\N�����*B�81��tI�|�)�U�ֵ�M~�t�Y��/�"��,�����,Fx�D��9i��A�3�~�7�g�ش��u?e4�����߰���wV�5BOto���:s��)H;��K���-_V�y�Of�v�؍�Dpݬ	�6|b=z9�a����c]��G�Rg�z���kĴ�܏t�d�'R�M��v�*EZ��~����1s<�k�)�6ոNE��fh�5�	��T�;�*�X����U��BA��D�0��q�����;twF7=|�:_��X����1����܂�%���x[��iy�w���x�	�R纙-������K����E#���I
���?ᜡՂ�z�T�<�v���"��1���l�ulw�3�F&.����������>�bГ51�,y5S9|�����ŉE��c�&ٍ��T�n��R�i�+��[8̇T1e9z�%׽!F�E�Z�	��&��x C&6�&cӦ�s�,gǖ��FX��sOq+.3��.vuP��\��$����"�g�+	0`��:�V!�2ݱn�5����3t�!��v ��,_96j��Ek��wZ9��솈�1�,xyqܢ�㻗L����I�
�o�?�����
���+�*�ŗjB�>dH�g+���~.	�(�c<����F洣�fRLJZ �=py}�Lw�Ķ$M�$�1�H��Oӱ`�_�<��U�J� !�I K��8�� �V��=�����Sw+}�I1YHѡVR%z�N��@yp�����h-�x�D)p>�#H�gڠihh�-�n�v�U���9�#J��´HZ��eУ�ŷ����m. ��zCg�-��Ǫ]㈅8M�:PĶ�_^�]�k������D�"�&,�!|!�$�z ����!��y�G�|(GW�ӕNe4�	��B�� +�Z�_����&h��8�FIs��_�;�����L�9���Z{�+56J&��k g��gJ�F��a���`z O4Q 1[�E�3��A!V���^� �V<��ҭŷ��y�3�._ɜq�J�~i�����:�%zEz����я�rS��##А=�U_��Qq.;@S����]/qDs���ۼ�N��F9 M?�1��~�����9ٕ��K���7M�@�T���"|�\�Z$� ��������
�_(���կ���jz�l1c�]�'��u�����U�������=i���h�{8W�Y:� B#vP嫛O5ǈB��$�y��s-��#�zm�A�ztZ4�:��t��`;T>�������C�\zzG�SX;�C�ݪΨW�}��0ّ��p,�1?���� �r�gB�q���U�le�����:��X)͹Q�#h�)S�Y�vQ�-����x %�f��*��b���l]T]D2p������g��$��V�}ϼD�Aʋ��})��6��92�_G���
���Xo쁾����w������Au��g��l���'6|\CX���2��}�c�܅�
7!f����5l����C��B)N��`��`�#�:�JV=6���U�ں%�N|��kz;a�崯g�/s{�v}Xk fa��|�R%xĬ�q��\��Qg!`��y�ON�j���u�$�a���)���d���B!"�Ʈ��`�X�OEM{�nw�!}N�'���łh�Q�(��Yv��	�j���_��r�]Ϳ���e9����>�"9K�b'5]�Z�_��;ŉGx�|3��4��!��с�C�����a[O�� ����n����&S�@�_���Ď�<�`�����Ʃv�3�/���4	�c��Ba�-���C��^8��	������{D�6�e:N!~K�8L��eM/Ƌ%�ѯ���)� n�r��T�x��U"4��@���×qF�,����5pZՠ�Hn��gI>[�@��}q�����yl������e�<�*�l$MZ�1���o'J��P����Ҝ{oM��HT"��:�F�ϟ�փ�#,�w����B�M��U��;��YQ"����Ě�kR6H?���:;D��8���q	H��ٮ�?��%� ;	s��L��A�� wS���<!{�y�|��>�a�"�Z�n���悼�0'_�o ��]6˔��Ī����*B���3A��uMc�^�d��Y +��;�G��G3g!�c�5�m�7�f5\U��૞;i�~��Чq���E���_�ca���p�(�J��^�9A_i��C<��W��ƺ�_�(4�{�J�'�g�J
+oԃ���8(��h�`/��XH?~�,�,+��	J,c u��?�-���d�K�lc�b�����E�R���_J9�m%2l�3lC}�M��hs�P�t���4�5qH�����),X�E���HP�����Q�V������WÑ2�M%������Xb@��l�6�I���p�l�b��Zd�n����=��Uoy��0���Um��v�Ձ�X~^�]�d|9beNTig���i�Uĉ+�p�FK
bX<$�~��u�#,�98��d�?�nI������,u~�l���2�5�]'O��#?��h)]�����t�����eS�e�T(���� ���l�e�S�>;L,�D�DOp���g�[Z���@$;�O��L�$;O?�n�x�8.�J��<��$؇������o'/n|S7�Զ-F�xr�&,�	�iv�o��7s$<S*��M��&�τM|��0�u��n���eL8���j����_?��VϦs��Q��$���eBI�9�o����e�F�ye��O��'#�*��Q#sd9�
Q��ʦ�¬�\]1����Wf�#핍�֟(�a���}$:)wG��	;K��(�U�6%H8a��fFd-Vu<�H���R����#��ę=��؟����^SJ%������&��o�Tvč ,[0��h�~�FӘ���N1ke����Gd�|w���2�z���R�����Ϟ�1.sR�ns���l9��Df���J~͂�V��[��K��W�S�PQ��1P��m��=p|�,��O�WR�/MJK����e(2A3�ܝh�vKB���˷z�����cf��-;�~�c��cיr��Rca5!������n��u��)�E��~���9�>54 ���=)K��?p��96�������6�AlXjnZ��kY;� �!��O*�����}x���/�x�1-�:�&>i�Q��(F$����˞'AG���`Xq]%�m�ɿÂ�Hȟ:d&0v�5kB������m�k�®�0�U�������랎>6�~���|�ڹ:��t}�4u��^�y����l�D01����G$;�@PBR⋑���@b���ݲy̑��&4�z�>2aZl����
���wH��7o�S����mOEf�Ьaz��S�ӿ��
m�6d�(��+�6Ve�����t�A�A���	|x>c5�?��䧐�&
�J���钞�:�}XŪr$�-:�t�� 0�:�|�;�9v�3�_gc�?ԏ+8�w�_�b�y}����>S�|t���>�HԠ����A/����Op��~#� �_�qj������ �;�<��x`��?�zV�p��b}����ƭ��J�m	�"��i(��xl��$�[���Z,��٢Jyk���k�* [�=GV��1_��=���}8�e�6��p�����'�5I��1HA?�$���)���Kʘ�P�!�QN*��:�]���|
q!��qU(SX�2>��W�C�]�E@R����4�^Ģ��7O�m��t�|	>���+�|�7T\O�et�'���ƪoL4~kl"	�?�&;��¯B����c����`ό��5.�p����XDm#tᰊ�VNR8����iL��{��r!2 ��'![�6t�'J�f�K$���ΚR�'�sU�Ǌ.y������9,��j�|8�Ln!�ݞ<ު�q��j	��Z瀾�ϯ�f�EH�D��DɄ��z�2���yYJ�����ʁH��e�ev�.-÷Lc�%]0�4�ߜ��A�������,\v�FB#a%�_j��Sփ��B$�_QgՇ��V����%��n�0r(�$$���Vk��Y�}ͥ��>k9��������c� D�m {֞�m|��V��*^8���j���,
`��j_���&�ϴD|�# r�e+
3���[��r���._Mjm�Z��_�HЎwuD� Dأ�~�"Ǩ�f��y�=Qy��5�0�o:���2n.b�Vhl��_� ��r�6ه����g�)N͡,C�6`���O��Z�o�	��X�>���=x�x����Ԕ,R��uQag�χ�����q�V�o����7��qiGG�f!�����[�����pE���C(���]�]���o*TOΥ��T;��>�˹F�Ѐ�(B7@Z���TD��
�o9�H���-Q.r�+�HSfJ�8�1+ߟ$��d⯛$�O��|8◡�ȗ�	�rV�N�
4�1T���ǈ�J2=�v:�TD����?8�G�<}Tu � �y��O�)��d��ݔ��`�Yp@�K���E�+��z�.�5o���e��;�v����E�y�3�mLL�ՄD�\>E��ym���	~&��kK���B�sx�d�z%cD�Mޙ����S��"�Y�H��)/8�d$��q����d�]T��*{����K�ӫC��HB�t5��L~,|ݍ�[ߩ�u�m����I���50�&����ᱮ�9�7y\�����{6~TM��H^�|��-�����}�A��#�r�k�\	��IϮ����"���[rP5p�a��M�A�`����(!�2�o�QQ� ��FLܷF�k%$a?W�c�̾<��!#�[>.P;�2z/���j7��J1��Q��t�S=����tC^��?��K �LP#�Ji�h���{�|q�p�]�E�w�<vNF�W�$��v����,�iv�ߌ��S����)�o�(��ؤ<���l5h-������G�%x���KǮ�.�%�~�@|l튔�:���@y�Tiv�膚sQ�mlr �NPv_3�}�j��.]R+'O�����@b+��`�`�H�;O�*�ѺW�y��&���jO��I�_}�����Eh��5S�пq[:v���i��Y��Oi�ߦ�lD����/ص/������L/��*���xB�n�T_�U��Qqͯ�������/w��`��gW�Il���Dw�t��_u�
��L���YW��T�hՅF��Y(xu,����k/�D��!A{JE_ʌ���:�����qzaT����kł݉�KM:�Rv��u�԰�lN:���.Ɠ���i�P=\+Y#{V����~��z̚�[��7����	��n�8R>d�3��Ԑ�`:�R��7KeHF��r@c\#�PD�J���n��|������L��A@����o�����޿Z�^�"]ߥ枺�������� �bf97��	��r e��%�o��|1BĲ�n�����]G���ϔ�v	�Ro����zv	L��"�n�*����ς���ىB4�����Ƙv��I�����'�t�]��e連	��i�^YG�mĽN�)�u�v�����������Q�����^���K�]�2v�D%�I]"��|A�p�+OK:QB�o��9#����?|������\ȁ��*�5Xy������҃�:��@�PJSyG�n@�̦/�uݽ����#:2��Qs��G��/tǾS�5����K�,�5/2��s��0N�%[�1r�2m��\Cd� ��NH�(� �:�ǲy��J�t��^K#�\N\��ꐲ�LGڍI(�R(�����7��s�˩y��zG&0�Ս⏹� }�S��E%.Υ�\��o����xA����f�a��c��U�j��+s1?'7�}1?բ�)W��><m|�ax煞� j�5�mF܎��N5�_CfJ
ER���������ګ��8~���A���y�V��V��H�z}'��wP����=���a�W<�Q�/M!������W���gȵU�e�h��HL��B{�&�t�H>��\1@��N�`h�!��h��q���a�)b���#�I�\9JpH�z(��>���"���KQXxo#Ԯj�JS/V��������m��I漮Z.b�Ѱ�?	X���O�,�o2m�����;,,���=�,�\9�׆����[� ]��7 W</¹��6����u������y6��8�X�e`����4���^�?��q��ݵ�?�aNK&Ӏ�$:H� ��=5�9��� ��DuNd�#��-�?!,k���I����\�pRե���(\�)����O��#Oڴ%.���<��Ox�H ����|�V[yI�IkU8��Gh�U`��ơ��X^��l�i~�����2�v��]���Y���r����:�:�9�/L����j(w>Ǩ�;I�a����5��K���Xe����|����?��i�9��E����]5S�RX����"*�'f�j�F�a��SaF�� ��E8�J����KmfƧ�"�P㓉���_%3"�(�8#�)�:��
�c294>O�e���T��`c	��BѸn�1T@k	�nȷkA�s85�lfP�tv����o,���oR�E��{mL��f��UX�K�_ʿ@��Q^���(��	��9y�+�Xݬ���EWW"��Sc�D��"' �;�_p����>��'%eL7�t}�d�{�Mk�@E����s*ȝ�n��GGzl�:�+�����!��ȝ�e�-���&�;S��ʫ�Q�;x��,�E�\�y��ֽ�oCF�(�1�`GA76W���Z�:�Yx�ugX�0���}�[��	�ۗ�,��� x�ey WCX�������o׃ng:�WHqxېF�YtY�"{�|�\��h�E��BF1z�E�UWz�wʅ����Nӈɗ �ݾG�S�+Y������3��󇥓�Q��ƍ���	��b��k7 `L��:m�\<��6���P9\���)Yq��8`C�~�/�<��~kJ4<Xd�!�96�-������~��	'�@��"�$|���7d��e3�5E� �*^���r���������)�K��0�w�~:�\�h8=�'�ut�N�~�f�,��s�:ÔV��S�i��w���8��b��0*���#�[���-u�W?E"��~�fɥ��~�I���Ήc�l�����I;��--H�L4љl�vt� ���V��[��Q�)�>����oҞ`W�8�����k�>�/�K� �,��2��H�f��[�.��*NtK*.9j( O�;~'ؚLg�gmΕ���b,l"f�]nW-��
JH���m�f��=̲C~n�Psq�pLCA�3d>�0Ç�/�wFw���c����m�d�<��p�/0���st����{)��St�a��+;zgN�ɏ�)��l�%��u�}V��yH޷K��&��2X��A�l}�&H�sP��$d�~�˘wW��^�~U�hm*�"���^+}^����b%��}�δ[%���Clm��À�ͤU�a�6�8Y�*τ5$���]ҹ�i������,�ov�C�8AC&�QQh������x�J=M��T+�,C?^�dF��&5�fe�I��3GP�O1��S�Y6���ʲ\{T{8��I����|���K'i��GQ��MB�!y�z���9��)ā�1F�i�����d�3�K}��g�!6?xM��mXB�UChL�s���7M��0п�v|�!���v �e���\)mA�|���K����ߴ���"s�EfE1y�}���q��o2�?�HN�,����I��K��&�,4n؆ �!�W�f��#����v�����ӍA����<[{�pJ���ԲS����V���vG�[8]��Lp A��)|42/����6#� ߸��o�?��(Lވ����������/�׼��=q;���'K'@C���f��0&?�T��\=����oG'��������H�JJ=�؁.�gA5���S� ��˸`���KaՀ�"Y�"�C(���t4�~��y<��pR4���32��:+��1 -e{���+�4	F\p����b�X���@��;�(�вMި�l��O�|l�~X�i��"���0^1�t嶫A�pSF����ſ�2y�?%zl�:�(�
v�Lr�K���^ڽ��R�$��J}ISE�P�GeX���X�����#��˴!c�Q��d
l-��xKN��*p"�>r.�t�S͝�N^�z-��5���V�\U��v��8ߏ���ݦQF��].��#��s!��ZZ�&���l^x^�����3���Oa@����8�M�����@��<v?,(���
��:��\��1��X�ݱ��|�ݫ�Bϡ�s�����Y0.��m�&i��}������O�'����]Z�ҕ6X|��E�����yA��]����3�"6"��|t���W�Q�����_>�L]_K���o�f�	�K�%�R��	�J-��G��(��^���~V7_Nd��0&OS"��BTɅF�VW�s^�#+z!P��i�Z�<��@�iݔ �g��箟�@�+���	��{5������Ag�p3�QN��a�8�Viy�C8�n h�d6���p*nS�u�|w�Ey*n'�Q��	�s6C�+N����#���ܰ�
�SN-Jk*H�OM��K�� ��~8Ʌe��^��r��$�����4����B�n�����]��n��3�z�a|�.7�)� ���V�hH
�]I�������H������8L�`6.*�5w�mҵg.�$��%�q�����JҎƬ�C+Z������q�O.���j���}�%j��D4J}��oY���1�j�aN�����+�]V1�`�W�`4�
���4�Q$��sDP��Gum���k>�
�K�]��Y����
}�X@<�-0�Ǭ��h�wuK �PVC�s��V��QP����:Q� Z$>'���C����n�͔��obP�W�~mt�|&�U��IȨC��nM��(�v�z��_h�8D��c֤�t���6�=�_�Zy�E8~s�Q.q���A��t�V�uM�b�࿞�i��?���r��՗��P@���s���8��,rEH$�i�BT=v�E-��+�h-`+&�G%��5�@:��WTwo+��Ӗsy�G�$�&EW`�kx�
-�`������̆X �*�m��(���$:?\�2�?���6��`ɖb�q���7Mͱ�'�-p�F��$'3�◍�B��P���,���usŢ���'�Q�pzWŲ|�|�o�% Ҝ}@/˿1����4�z�!��ٱq���{��8ԉ� ������.#�	��ԈR��eĽ���X=�eCϝ�mUG5FM��ێӬi�-8?|�	�Wr��+����|�\�������1����"�PӯJ��eQ_
�S���!�n��ph�xA@6�y�8^�o��\	h��D�B$7�y��G ��S4��6��`Ө/�sΗd��o9���!P5�֑�`!0�$H����:ƙƭ��Mԙ�s��U�.]�*�3|��:ڠy��5�p�K���Z�CO��	^��:���O��nݸ��sö́�[ԇH���GB����#mw�n�<�Dv^�9}�cE-��P���U�O�6/������nGM��"���<�l67�y.���N��B��qfh.��d�cmEހ��g�l��;��|�O%��`�)<	��E��)�W�C�jhe"�������W��L����?d+�B�]�NI�X��C�B9;�����j$4�S�d��969w-
�G�W���\G��<]���1%&�vX��&C'��3���������ă��#�lT-E`O)�o?��eA�)�X�5��?��n�8�-ds	kg�����4I3��<B|����r"�._ý	^N9,7o:_��UF�H)a��b �蓴�mG:����Ł�P^S��]n7a��:W�D�	i7�s	���X����^�G��9{�=Nz��M<YY�!�J��mv��)�����t����I5*��rVsT6zY�S15Rx=�̱�t�3xQG� �������M+�Y�VL5�?���5���.ZT	���n?\��5KV��C�������с��%
=�6/9�E��6)h�ہ��`��v2��o3D��~�G�����A"�wH3?9au?�_A��g�c��u��:�q�풾=T���xt)��Ɛ��0[6����>�
#lٙ���{��Fɓ'��V�&ד�#�� [Q��AtkT/���{�U�e�(��l7u�n��<΋�����"ӪX�����F�$P$Շ�Z�p�F,JI��20�����H�/�J�>����̾�� �n�)�:+B�s�4���������/;?���b��O]���x���g��R�-��2֡@h�8ь_l�+��K:8(wg��AȔ\��4m������yǢ�%<\jx��݇)qhq�.yF�l:[ 4�?W�'��8	�N�|\Ѥ�k�?���: ց��.<�E`�d�IJª�Z¨/B<�>�T*�����El*؛Dd_A�1敼H��Ɋ%6OAW��S�+��;�B�|�ܔ1�ߓ��Ԁ�w���ϔ8��f�ڼ��d��E3�N���*�#T��y�j? dW0%���� �u�ю�SM�\���� :N�j���d�LP_���[M�2�qZ���M*��"uju�(I��7�=BEM������e���M��NR0GfкGx� �VX�ٗ���7�������F!/Ŗ�o�w��;�@��U�ِ�ɳe����ul�=;��;�X�.g��������cj�(]�"�	��KcE�B�0� z�DTqĀ������o0��s��ٰP��+-����R8|�D:���2��K]�x��[��6�jm��>������r��n�Ѕ;
�J��»���!�lv�H+}����D����u@���um|�֨� _#(�qע�Zf�d%ae#�wrr��2��̹�=�0Kx}6g�i��K��� +.�fb�q�K�N1�6�:y��2����-�5�X"ppJ�u���Zˊ�Zx��r؊�=�-08���.xP�{�&[!܅�d���]~$�%�m6wv��;������\T�������&$.~�Iԥ�� �9�S>��ja��ƵI��݉�ͥ:��M��/*ϒ��#B�ӊ+�<�'V��"�/�ܜٗ/��o��i�]�B�Rv�R�UN.sk:��Kj��Ef��c-w���arTu�T;Sr�A@���H�b��� �X�h��\��o1D�n�����^;� �z��5�A���u.p�L2;/`���WJ�4�W4~;6����.e|��`��s��5�}�2'�@'0W�H�h�|t�O��;�b�T��� �SW�9�����7�	2�x>OM�v�I��g�$Û�2r��T���(���%_ ��>�=fG�W&N1,�k�ϓ��	(�\y�n%-��>���Wg8��S)�E R)���ɞ5�b�	���pr.c�7�!���H��^K���__�.�y��	�^^%� G���:�� {�Ua|�I}^�V ;Sρ�\�$ހ�����]FG}�/QQ�֙�r�G�[���̾a�Uk�=�0y�� ��z�~���HFE�̶��컿�qa��;��K��=^MTޛ|���ۭZ��쇑�S�鸁����Q9�Xx����C��/ӂ���ڻ��v�S4��e
7�Y����1۩j�k'�vjX��n�K��-�[g	����V�Al�t���	�Ei*qLM�w��N�J�;=m��۩r���6�X����X�ҥz& ���֡��v&RG��M6�JgR�s� �4��v��Vk�-�ۥ:�WysV��LE5�Q
6��n�m�ŭ`H�d��@���i��}�#k�?��xEpמw�ƚ.`�a�J)�4�Y[)_|ِ�T�C��������]��Pt�8p	�\H�X���&�gG
�PN#���l>�U��b�/��\=Z�v��NK�k�K�|5��P4=[�XE7(�
ll#�CP��2��$����D(�����a�H�<}*�K'���쯴I�퀓�c�h]*QF�#Ld���]�B	/�U���3��q�xz�x�[?´�~?ˈ���R��X�J`7�!
gR�o���R�\dF4V���ܾ���PX�R�~�:C/�+�H�T��Fy�&�(���l�y������Y`Y��x��l�_���B&6�^ �+¤�'��డ��(���;/{C�k�v� �D�l'�V)A���z�U�CM��Ґܻ���=\F;-��N[���Ƚ���6�%R��?�s���*:l���Y;ez�*E�؝�O>�ϭ�r�3���E���G;TM�S/NVBo��s��Wj���K��f����ǾC�Nl-7bi4Gù2��#@ �k��Fm,�lH�	V��$�	��S���amO��7�M�ƲS��h��S}fͯвE���NZiv� ���
(�cg��{E���$��k���{�?\G;C>��v3����� ȖF��ߕ�������\�L?�Av�;pk���B�盠�q�T��K���sn�yn��
ʊi&E������k������@��c�x�ߓݴ�����O&uc��cT,Ĳ��i\��B�y�B�y��׊�v\��[���k]{�4��
>�c��u1�n��k�˿2��C4��qh�+h�Ӈ_��^ނ�QG�Ϙb����J3YIq-�Q��	\ҕ��s�w�D��D���Ô�cqԦZR��!N|9�ݟXT�0r#��� (�S{x��VٺJ݂�yU���o[�6������d�Y#x�%�� �3��9����5B�G��ۣ<�#|����q1�[�Y�����F������"�<�Jm���3�د{)Ғ��5�D�?782�DU�j@��%!���/�!�wpx�n�[�N4��6f�.�pa����L%h��-�5e�δ�~��Oq_9�������9k'qC^�q�Z�Z�6^��І��=���$m!��>�av��!�� A�k!v	����p����/�pi��=q�S��D��Y��Y��ma3ʡ\?RSb�� ���^��N�>�yo�*VST��<��v=�JO�n9�X(T��U�s���{�5���L�G�k�,��?��n�<�y)�'W�R��x�ðsk`wf� Y[x޷�`�hi�S�8�#��CC�y��R+x�ϭ(�x�{s]�ܐ��V�E���9)%;�f�t��+$Md\�U���ܤP���WZ��ˣM{5^q��nG�8=��I��|<��H}��A\(i֪N$<t͑��P~�RR�q�J]P&�5+.�^��(����N`�����ӟ<c�'��G��>�*���Zg�W�+�_C��{�ب�M�ͫy0��B��� B(ig�����wֳi�b;�t�,|APw51;�Ӂ���a��o�N;�ol��`)7Hp���W���>�>���-5u%�
�����{���'i��6�kb�g"B�����?� �\kM�-��`\��U
_$+��=�0P�̈́�Vr��Ë��X��0�������2r����e�:<,�/�5ST�6�1�H���S.�!��3$��Q��۹�h0#N{(���SBw�gק3҇Rmp ��\	3$���r�ޝ����oB�v�6��x�[%��:�l��ď���f��(9��KS	L9��p �(+�<1�|���~>I&ZvZ��s��F���T��$��[.(f�xTЀ)Z���x���#V�`U��\�o"�����!� Lw#E�	�b�IM��ȩ�����X xq=�sw�1C��
h������W]L{�-$�F��d��os�R����p�f���=�2w�n�}3�6��Z�g�`s�Z����N� D0����%���x�����:�F�J�����W���}���T��'�<���|����P�5I?p
���bw�p�Ⱥ@�s1��v�%����L�]濔��w �2J�� n;
q�"��{���s����Z,�@�w���	��s+^��C��eb��ߒ�5Z�ˡ��v��k���#��
M&����,���y�\���f`1Ԅ��u�Z��O�
������N�C�c�
g=!�?�
F $�H&��R�E�+�[F���ֆ�:q����~vFQ�ϾjU��u��� 96f�d��{7C����������KSW���3��s��#�uװ�8�J3���i ��G�`R!�5��a���hhK�ԧ�<9c}�[� QG�Ԣ��y�A�ɿ@1ߜ�L��q]p��y�Z']�[�gp��V�ӒK٢u���J Y���V39`{j[r�6N��T���[r�c��g{�"��'(Ȇ+@���2(o�E��J@1Z���[�Y� A@�^�ݨ0����c��]]^D��i���O��:7n,;}��[���bA�c0O�z
iS����cH>�0��ԡ�m%H3�x�{9E�5+XQ��@��@_F�"���F�3���P�{M�l�Q�w[�d),���6B�����~U���j���pr@��˦�BwZ�}�C��� 2�w����ʭ��$�||���[�hwN��� �d>t�V,)亐[��uA�WM�~��$a[4���T��[oݶ�v
��QE�6��+ 0��"�x;�ȍ9Sn�r`�|�D@�D�������č0���*���.��e^�]����N�L�3p��1��6�AtAC�/��f�<�Nti�K9���s�< �<�6�L��������M�yW�������Y��TZ�b~f49��=xi˵�(C�_�� Q>���Y�A����6��	�A��敽8�0K��(�w�W��O��h�'�}��8D*/v��4����
E�xÝ?���Z� �m�&5?��m��O�+ͅ��Zl�,���.�E�4	%LN(��$f�wiP$Ҭ"���0ȋ�����?�����T����t�����@b�^1�_/�o> I�ғ�����~�v�K������lS�u���7盋\i1ͳ�ȺW�"  kz@|�a.�1�E��UkN���;�(MY�`czz���'Q�9�[+~�|�,h9��*��V�P�y�y�؋�?{Z��R7#�T�O��8����,F��\����)�B�b�	K����rB G�(�3������&k�(�p�/MbS^�B��-�p���L�ǩ,~	8�@Sw�&W�1�Ȭ�_og��%0Xx���w1�R}9�AO���;�A�*|1�܃�X&fb2`S@�mE���7�,�(�8K	"W6�ܚ�(���&^��<&�q)5<�r~�S\`%��V��.14�ޔ�q���WL���j�xH��cs�Nmq�#4����դ�Ƈ蟫L�����K��&nb���l-���'���)*Ţ04�<�GI6&��qX׉�O�Q� �*G�U��zt���)���Բ����Ӻ�HT����C���Zz��s#T{t�*�=6U��i`wqLs>��?���85�Vmj�r�"]�()R跲Yk<� c�g�1g�W���<�nZL��[�#Kī+#��FZ�$y��m}�q	\R����^B����q:����s��b���?����RO쥵FgZx�D����6HF��	���!��_n�PP�U��C.���y��@t��DC��ԑIf�/�̒A��I��NЅ�A�ɜ�� 8���Hxg�b4�j:#�����Im��T��gN�\Q�1�8S85����p���sߡi�ԭva��y��x�1��d��H�Z����x�|v�N �7]�7����飄���f�����I�y�6�ܖ���.��b���v��Q^��]��������-���i18z�ݚ�Zt��b�qj������,��LO����Xı�Y�c��N�����4����{�w/3���$��b5T��?�|H&�%��Ja�躾)���(MVsP�63�-/
_FTH� ���(U�gԜ6�ĉ�h�U)�5))oʼ�ʬ��C�o����vrT���E�$#�eQ�N%������P���R��z���U������Z�%���j^�����ʸr��i"'O$���Z�Yc5GG�s�bD5�7�y�< r'�%�X� k-�*�{�i݃�?�!��\~��@�x�d�Md���K�-f��1u 7������^?#�3lj����U�Bs�uy2�w��ׅ.ֹ�G�;PT�q�8M�A�N�z/YNT@˻g��݂cp2Nꢉ�0m�):�88� ���@Ҙ�?��b��ud"&-�X� v\�د0� 0'C-X������Ap�M0�2�E/x�VwP>��b�3Y�~�!*�J��m^NN۫�w�w��<\2�RLM�fj�8.��D�3�Ҙ��w�m�bmg�2�b\Hmġ�\�Z��w������������OT'
k�4��)�"�^x�ߋU�u��x�6D��qt�SO��J4�Jo	�-_�L���4��n9Wܿ�a^�+8RQ�r��vn��ҍW�:�+�MYS�Am��^}b]s�j��=-Ȃn���;*Q&�KT{������Fx��;�}m���ޅ�=���� ӃNC��S�v��c]1���[�r
N��,�����y���I@�_�C!h�V*�T��:s�D�f�AIC��d:vo�:��嚿C� K�甃�奶f�b����e�̨�����۵z9-l���UH�/N�$'�T���)(��ٷ�5E�Մ6Wr���k,Ƌ���k�Շ�>��~�*'���n(3��!#�Y��� �Ad9�,*�F�0���:-ig$:�Z�2��̵��⥮T�7���G�޷4�L�&�@DZ�g�c�7�� �3ʹN�ջM�Γ�J~���� Gn��"������t�G���N�b�N��F�G��E�gc�S��$�M�e^q1�X�t��e�I�����:�t�Ϳ�:n�P�?e�VB�6�c�&K��GC2�|]�e�]� Z|)N�&�3R��Q���k.XE!�d�h'E`t���*y 0�) ۵J���r�u�R��_�M��u8�c[����њ|��Ӝ��9�)�7]�1�p�;"��O�
 ���
��B���'.J �dо����Y2l=�;+�+�-�
���<�=�LRc.�h�1`�=�'�����4
�x��`��2�@�k�/�#���S�0�-�NR�(na�Z>��p��Y�͵��G&$E�$��~j��[��������AȸڨV{�#��yޝ�G\�U���[��.b�T��<�)�FF=��{��84 �N�@=G���d�
�O�f���L�p<^���cP< �)ɉ)0f.��l��Jd�i�Ol�@�zqI$���9p��f=%��SͰ��YŒ�3�3�<�a��P¤�P�Gx��	؇�_��<�.��0e���S�mD��V�qv����r	p���U0�X�lV�:�( o@�������۵4����g�����	��1OIW^��pn��~��~D� 0T3�����G;��Ř��|��Ή:�ë~mSME�"2BB@q�j�B�}#��8�L�� �IZ��/^b�#��f]E	�����.0Y2´�*(uq�1+j?����i�c���*��]B'=q=юI��C����ɘ/�B��F�7�fx^VVL����0�3|:t5�����z��^O��2;iIe
��h�?�4x���*Rbo�p-�uO�����?n+����o�_Q����U��0t��ۏ�u"�x�͡_��Yզ[X�E��� ��8����%� ��%.�t�W��樑�jְA}�ڧ1��!��
�z�c�Oⱻ![����A�������PW=�Gc�j���.｡��G,��%z1��A����G|�
	�9�J�z)� 2#�M�P�~A��)-��ţ����]�e[j*	I{2�lp[BS�<����r�'�'i%�:��1��c�+J��o���F�p�x�Vn�S7n�� 6a����.k4��Ԑ��Wb@���0�����ͧ�6��
>Ŗ���'T�q���+�����Ԙ�+��DL��h��Vd��4=�n�ד�Z"F�����.�J�Aӽ(Ml{�� �;��2:nl7������o)a����@��3X�㡏R�L�T�_�V���������P2��IUFk�<�*o�1��w��>���(�5o��P���:�a�H�4��MO���'� 0��}	��p}��& `��[�M1d���T��W�����f{g"�S���%��I�mV9�2�B��`D�� ��'�����=o;k�F��7��%V�ؓ�Z)���w��@��h��k��&{��K�|�!a�u �����>����&��b�$��u1���"<�Ft���Q���C7Ky�Q�i�^����(�j��i��I�A���3���A�oK�\~e�!,���w�e���!��r�������m�F	eI�H�0����e�b:��]�`��R�\�����>/�l�mr�z���L�h1NiS!/X��[��0�\��)��z��8c��`tIO�.�7��/�!c��B�R�Ȁ��w=("��uf8�5_��e����O���t���+`�%Kac����@ei+��Pvܱ��K����Y|���r7���;�f(+���/cWz���]�
��Q�0(VT�����sq��W1�+�>�zƂoPw�3��lc���'x�0�Ԟ�����z�/�^�ѵ1������\?_�k�o#���>x�w���m�H��9?�X[a=���*�|�b���G3gC���E��s���ԥ����/�������td8��-jC���h֫��&pJ����6K�JgX^z�ym��)���ث}�����ȴc�|�7:��R��"W9)�v�f����%3����Q2a��ʓO��/"��nrR9g�Q����A�A�B%�Π)�p<
V��ed��,�z�s������.\��"�,�G�l=��V���H�z�vJO�ͬa��WӺ9]h��a�E���%!���7�O@�����+�� K(���]��g6ﯿ���}ʗ���lt�w���C_���4φzW���3������?�N��d��\����4�p��h����>��a�[]�}�pJ�ՖL�>���Ǭl�}������#��R$���B��<�hQ���AD� �eЪ�[��e^HE�����(�}:%�^v��C �8�W�%��
�Vs�H.?�N���@XWU��a��o?�e���%�놔�~�뛚#�z~���w���
��.In⎐�P;�T�	�^<pZ`��t\sL��韷{U �S�$n���zJa�%T��Ǯ}�WK��#̤5Gc����@y����Q���Ca���w��k��3Q��Ǹ����Hr����0*�G�Ö�IP	�IdT�/}�a
�(l��ps:N��2h�����S���j�P{�5�>S��/}.`U��ߓ���$������O���(z
�R�AT�-9HP��(r@��66��y�Y2w��M�[��u��kћ��)?�׼�'y��/�dɥP4�|3�&xrҜ˶LYq*1��_��T�:o���n�Ic���6R�NW��Xh��N�V�<���z�XB��l��j��O�}��@��_��&?��3W��lk�Z���5�ޚ�
�o���;�hwN�VK�m��s�x��ڠ��7�z��'S���͍G��9jWC��G���Kf�%MX�*���h��n74��\k���M��0��Mi�D��j�����=8�h#)�U��c�����Y%��@'��s����0�ʣ�Y��?#�+�T�{�*{�J6�7�-A!�ܥ����lS���b�:�Y���T�I�t�{4-=a�%�z�ʩ�����C�EN�>����]1�����>���r��Q�i}+qP�r��{�Ɉ<8#�9>�s�[w�iL ]���&fQQF҉x��┩6�M����A�Q�'.v�?gd��Y��2�1��뷳T��Éجn�	x i�ٷf����ߗr���M���h���lI�ד��C��H(�)~����{,G��-����H؄��q�۹M�Z{Tu��*xᛂ	��zӻ�|o�p�ʓ����鸿�p�z�)�l� '9��@i<.L]�}�hx#մ���	> �"�~8�O��d�qԡ ٮ*��e�&C��^'#:>�'ݿ�^d�єN+A+p������e�g��]�>��i�L�D�Q�S��1��ϣC��b�rb��s�Ɉ쫭�0��C���mq�f�����8F�m��}�^7	�_�ES��l���s�	�����<���Ek�GД�F=P��Y�y���EWm�B�z�2��z�vG#P\l����1VZ��v�h��U�)���G�Մ��� ��;�����.wԙ���[ҟ��l �Ebȟ$)���(kn��U7�x!x��J8�*�H����B�b�N�̟�r����zj&d�ψ?��4tC��šт�mn�\��l��I�3jV5�k�!��)e����� ���;o�/��Q!��y �]�r1�yx��B�/ ;<j�������т?!o��"(��|�;�+�?��D8fes��#��7F��ӱ=X|��.�g�o����<Jq�[
J���w��;�g.��Q��z�K��P���|������߬+�+O��<������y����(m9���Q�b���P�߉�c{�,�1�v섂-��H~ۼ����1��X#�M��4�"�"5�	dvZ�3�����(�[�c�6��v�z1g�|;J[�$�"�7_(��N� ���ȁ���߂ڲ�l&���~����խ�fn�m�)1M�M��������#�� C.�N����c-�rz�6�ʷ�I�Q��˪��";=������:[n�B��z$�x)�����J�TCw���R�{��d[jcCi:�\+t�o�~�N��s��\�Y�_-�Z��"
G�)��� ���,dCɾS���8h�t����\�G��ю�G�+��C�<
d�f�u*�d�j�'��W0���Չ*%�;�8upk�,�?3]��CI�0�!�C�Y����[3�cڟN�������`-����|P{�E�W�X1�i��%� �k!"��u�%�?$�c����d�߾0�ꨥ�spNK�.��$��N��2bq�2+4q���#*I���&�PJJ���%g�='k���	���Y|�q�X�V���n$�z�h9��d����$A]��}a�g\Z[".٪�og�����F��S� {�.r��X��b���A���)��������협C`O+� �O�a
\�VÊ�qF4s�p�*�w������3ţT��p(�U�!�P.LL����n�8iR9FьT�"�v�T�l\fR�U9@��Ԥ(�
<�)��M��]g��m����S �$:I���efil����#'7>������ ����]p�%|��_��wg>e_.��6!���5��J7�Nt�k�!W��sӹ��, 	a�*m��X�շ��UwYt�qb�+��)�2�R�t�Mk�����mkr�Ɛ}��M���?�NSc&|����bJr�ա�����K�X'9^��1�5t^�Hf �`���ܼ����Io��
YԆYd������T�1���'`h)]��}����x޷c��hp���d�Z2��W�� "m���G!��s�}�槈���r��},�':��%�Յz-��A�k.���_�aSa��{}�G\oRW�<�Y$��*�8�ey�����x�I��  ��J$�Ø�ÿo�C���4߇�����Jr��
(�h�1�r��KϬm-��?��~�cHx�%��k<n�&p�3�V�?6a
Y6{�L>��nMM
�jH�EDG��Rl�pzX�K��^�){��z5��ϴ�_��C���B��R�}ʮ�����b3�nI�(籟)5Ӽ2��e�v�?&J�dd��\���������������1#��.�Gۿϓ�@��_A;����֮��'�W9�U��DuI�S<_|oW�����"�;��/���َ�G��-�{��� ^>媃� ����R��\K�5��1���Cp�����g��`�˙�P�A�Fҫ�g���E����V���mH`}N�C*�nF`� ��C���T�2޷lV\�6�W�38�?rio����?����v��AK�"Թ%a��(����6�̪c�ѭ��i�1Iz����Sc�����Q�L�o�S��\JcA��ݘ8,>����Ҳ�Ć$��Cf��W̍A�M��y��D�2��YKF��ȋLV���X$M���VS�jC4�T~-O<SN��Y�/Rk���������YȰ8�v/�b-��-Q�W�G꘍0��O�(2�����%e�n�h:�¸��J����Ջ'�DZhTr����[��M/��.}���	����UM��/w����R����f�b�U���'1Mී�䄢]b� l0�hV�a~(ӗw��dT8D�P�b ���}G��7ز�U�3y�L�����d�R=y\Qwa�#�e�f�ֽG����@�Qs�n�B�u����
�*:yF?3�M&٠�ab	����9�?#z���~�%q��ѢdG�����D�(�T�+�G��_��Dz�7w�b3A]�}ۘ���N����M��֏?wC'ѓ�D	�K/���.�2���A��3��й�=��� 
�g�s�P9o�:g�P���?��
8�t%��b�zy0E���9����)��*�X�*+����c�OW %BK��fXN �cZ�d�Ya���C�{�<�J�d����Z��U9�x�B���|���Ph�PUm�</ \�	���p����Y�~%Hg1�=��xaA7E'
�ʐ�R�=b���OW�Tα?S(�t�g�B�  k֔¼ |S��pJfj��u:�q�Xva6��Ue����8,0z}s��2v8�1{>1T�ug������,�0&��Ĉ�p��P7�$�V.��	�[���Z���V�o�Ht+)�ϴ}���J���/��vnGAJ�:����Uu��G�9� X�T��;��9�o����#W��^7�K�a=Ӛ������-u꡴n�55 ���O*�^|�w�A��,61:���Y�Y�jκ��%9% v.M��Q�
�ى�?����e����x��o��;��R"�VB�@? �9�qĥ�<�Љ�K�Z�FJ���  _�Q"Ү%�y��a2/�pVs�P�eD��dè���R2 ���#�6B��5N�[��K�g,�W��fe�aB	;�C��H��wd*aC�p�2/A�������~��Q�Er�w��j��rT^DgX�\�!�5���\צhZ�]�fl<�S*���,U$kK�Csu��,�U�VT�%�RC5��JXy�2��%N�Ds�6aҚ�]�#A��!7oۙM��K�1�����3-~��?(Un?�:���.Nk����ln2�Ϸ��∵�4 rp~�NY��bT��<��[���i���NG����H���AX�D�2�IK(X�}r�!���Q�VL����Jk%���G���v�6 8�a��ޯ�D|o���aO~�$�v��r��!c+��|�n�k�iI<=�]��CdQ�t�uO9��#�ߛ�c��mi�N���Z��S��>�S"¯�U<�?�E����e2���*��� �`껿ϦF(	�C��B���
Vb�BLH�/���{��; OA�\��QH�$�z�e`�z�h�����M\����A�$�����q���Z5g鷳&�{m�ф��5u�r��ا��'�7�W�k�*vtv�0i!�(_̽�:Y ���r�3v�Sr���$�*�\vǆ�Xxǵ�� �^��ugJB�:Kw������S���x�Ųo61�(���
�=�()p0hd"@|P+?x���;��{��7��h`a�
As�-�0+��\��x�c������m�������5���b�[���u�g��D�N"2���ca�L����9��q�Ƕ1fK��?��>��+hR�����I8�]W� }�݆�3��m*��췽Ga`F�����n�]����R��q�m��e���}�ur9��wuvB��\]&x��O� wz_�{��2�AJ�
��a����lxkD�8�SE�~ի�<��g�����s4�f�@#48�iz�7�+���
�{�3�E��ȿ��k�GD�}���h�,��~L�͓:N?�j��eS9�*\8"O����U0�LVJ!�ҥ���j���f�?���?��_�d���r��C�x	����K_F�v�nM��`�}z��a��Y��8f؛��z̀J�E�H����g��=����q�`��ם2�qj&�_�6a�t� ;r�4���)��3�w"���(���6�<�T�K�Α�I���Ѓ7o+]Aҹ�����H��~50v��m�k�m�-��	�Q�"�<�j���z
,&��@t>���Y9�8 $��4�%�)y����t" �ft�x��n��Pl7�Ĝ.�ǫ���)��֦U����E�Y؈4F�C#�(��������e�6�L��2X��XU��ls$���|���jR�g0"
g�<���c2���0y����t�2�=�bA.��j62��L��Y�+�fC�aK�4��2�������!��X����U⵴��`�/()v:TwH�6u�o-�),��ﾯ�+	�;�b9-d��`KO���^{�!���Z~��3L�2Q�{�cZ��g�<����r�b���R\���y�'ޛ����7�����#�<��oh�j�W|��	�|FU�a�poF�!G�C7�C~�,v�>!u�c��������'��r"F3CaǕJ�;|@�w=#d]���%�TW/>���I��<S�4�N�i�Q���Fb��Ig��P��9F4B���F�+ ����&,p���tf�|�vZ�����f,�O�O%�CF�������*��$.4����z4;!���c@i�q�I��	�@�i9A�6G$���R�^�������Pv�Ɠ�}�+(����ō��@�ԝxy�;�DA�?����LU�Fc�^�?�왈w�]���n+�O�g��D��I%l�ԉo�����kڎ+B��t����q�f`"Uص2��[+�ַ�D_[���x�����W�{�L�}�`�����ỡO�{�5r����G �K~7���b��xc�Z��Ӏ��M5�桛��	#�g_��m���;�����W��{���2S�P�֣$��T⏾����>��Ʉ��5_,�lRAGťJ���Ha
�77S�3��M�ъB��������-�[�e>ˢ02���u���Pi$Hxg'U8%�̙T��O(}6�� ��gE_�HEy�m�J,%�`Ĺ�}�Z���	Lm`����xMc����=$[�d�G�>��9�'�$fI.	������n����<��f!�RX��v�&��rXEW��H�����7=u�GQ��N;�_�@Jkh-�wPE\Q=�gAs�:ʕY"h�d|��"�6�T��v'���4U��ƸZN٪���I~RӪCF�c�l�x�i�ZV�pZ
�d����!*��8��_mdSseI��ss�Q�,�Ťn�,�A�ހ�a\���p����o����mP�A\AW�wؙ�!zM����kj�(d��-�352���7e�'�u}���q�(���P�J��G�o�r���� ���xm3ݮ���6S�*Յ�3��5r�5�!;�!\ 邩�O�[�E�
��F�tx�6�<��n@\�E���Or2����ʡR�P�(���?Y�$��+������(�ɎW:�9G�HJ�r8��t�1g�XE��۬as��ő-.9��" ~��؇ԅ��n�R0�:��D@]̘-�0��>v�1�#�� `����ܪ��Qv_�r�.��adA����)�Ӏ����\^R;�|`�A�/8(����&�I���Q|�.�Ƞ?7?p�R{gǍ)R�ro��G&�x��3Lۺ��12~ˤ��ؤ>������3V�̴n��~��G�Р�6�5���!�׋�/���
�&���AE6A�{�li�8<�<_��c��-�^%8f��$�L��N��P��h%�	��'�B��aS
#�Ah)\n{�X;Hz6���TK��Yjn6��K�9�;,K�����ڴ;�"��������}�0Np��(������㍨*ɕ�d簸Ÿ��ľ�>��!��w��F��V��W��2�C�(���]�o���s��Ɇ�9������g�z��^O�_V���� ����yUdO�jEpi�'D���p�[j��\C*��[�F]���uZ��e	�9I��rwa`v~w�Y��t���;_�:7G|����=�m�J�@;5kp�s$ǀc��W&�)���+yA�{���^�j@����u�Pz�l�;Q�͟���,^7��M��E[@��vǸ�|)hϕ5+���-I���,�C�.ã���Ӫ*�C���Hl�Ʀ}�y�r�#:�$?��@�Jq�'.9w w=̻���p�}���y��ӱc��8Ρ�?֖I���[�7Ң�r1��i;����=�$����� ��(JC��\�l��q���U�	p5���F���� �'\�v"F��|rB���Z���Ý�_�� �Uߌ���zE%e��T,����xlQWf6�H�^!��/T�Tv�?���n�OExŵ5��c�a�Y�wM *���?��g��ѵsy���Ou��=��]�k�	%�[��c�M���Qv��e�!����E�K���a�өv�*A'o�k?��~K��P:�-�gq.˭&,Y[p��(3f��tw(��\��P�I���ep���9:e.���Tr�V��L�-�
�_	\JI�����Nm�W�<
�`�+cF�o	΁0j�6�0�;�;��="9����,=�\�֛�!I���Ve^���P3hSgl�^a|A��O��Ң2�XY(�:�>���Eb�r��L��O�)�"s�5�Ef��J ��$�Qˬ��3�b{���Ɖ�V7P���{���, m+����1L�9'ǵ�V0�e�hR&��E��Utv���^�Q�۬����?��"�	�o�x�U��f�F�f�:�˛�Lr�ESӨ �=hূ4e)p�YPs]����D?�%��Ȋ��m��aeJ�ZAd3v�%�S$���V�z�@�;�{��q1!)zM^�G��R�Y�J��YLL-�8$��͗�S��z"LA��T�A}!s���ڿ�$�m�,�^��'���=��p�:U����R~7�}��{2Ӂ�ɯD��I�+�Ն��oН����V�"�l@2�Y�k�5R��~eRlS%��AH��f�l��oT��?Jѥ����LAg�qʍ��1i�y����5��_�2u���-#4\]�W6��|�r�"��˶�\C�:����{�ߵ%j{X����J��m�x�8+��%x.\����� w����v��)J����/���1�$�\|g��Q�7�{5^�9r|�q�׃�kq�<�G�2�s�o6���
�T�� ���Il�1�����-�\b:�X�Y1��.�\tp�7~/_�p����,�j̵R��'�:�u�mI�r�tI��=�~���t\����'x��:`�u����:���X��!yK��@��C��T���FKu���Dn��$���s
�6�)�#���i��Ū_����h�)���'�J�C��� 冷��)�� ��[ X2��������N������_
�$���8q-�5�d�5M��~�;uW�0����>�r��Rک/�L���,Y�#���
�,YD����U���sS�"h�� �3��N��5Q����m8�O������Vi���z�	����+E����(`�}��"_��|eu�LZ��$ϫ2\[�]�<���f�~�.&<=6��f>��¶}�v��-�Z�U��&!��|��x�t+�
���
b��q�̍X��/�5��y�jgh#��B��o�s;l�_�r�f� qZ���B���U�k>'�y��F�<�GB���N����剝��ߝ����!�U|��zd1+i����+���s�f>L��೔����
�8#��Ʌ���!m�YQ b�rZI��� ���8��[�竂��!���l�f��kA�#��cўg���__Tꏕ�\$�=�����,�k1Ψ5�L���T��sZ�� ��H+D~�+�"���n���o7�	8pk�tk%2�'W��<*��I�!�&�_8l�*$�#ɾ��X�1�0 .S���{\=�3���%���e��@��f���U=�g�s�I�v�_%�iG�IC�yy���h��#�}C5o$\��T�om��M��լ�V���x��׭��0�'/���\��]�2ٜ%1]� ��BS��f�q]1!�R����z�2r��W��7	�s�m� s)R#�*�C-��U�����(X�$l�}l~�i��"\�Mਈ\O	C����*���uTq#<2�����?�rS���p���c����Q�
GAr_����Wv�9�S��m �j�^zԔ� ��n��c���&�L8<����r��o:)H��2���r<Z(<.�Is�:Ov�����f���

Ŋ����!OP|?k�ئ�Psw¯t`���R�탏$S���63���XX.�2a�N�"��Ǳ~�Sb=Nd����bW���#�'�kր�o�4;9H��+{��mS۩&vP�"�x�sE��f�������6�o�D��"����X�F�Xڅ(�����s�f�~�6�9�b=_�..h���ibL�� 7cY;�S�4?��8�Ip�#y�_;�в�L���٭'60O�$�T}��3
�[!���x�!��w��z�SNx���A��k�ǞI�X����r�KnyΓ�kE���1��
���:������L�*$dW�WS`� �%�]`����Y�¦�$�lztl����)�[Xp�,�$sm������L�C��E���6g쳒��A\(���)����#�Jz���b�P��"��1�xUC��B�� �i�9;�rm��+���4����P��х3�����2\"@�n���V0�/��5��r��l�
ex����U�}�.���V�q�3>ɆI����qmQ켛I. �;Ї%�K�j($�-̀����Z�g����_�^w��/g�@~��ݬ�*y�1��ہ�/���?�G��D`fy��q)�}r�0���t��%��P;8udtpY��S�4���q�/	w��rh'�	�H����	��눝}�Ra-� LHA��:���j� ���`&�fΚ����'�a	��#l���T�W�K*AHfb���X�?��85W3;(ٖ�q0l�r]cl��/�c%���^���+|��it_�I��S����n� h������qM�,oFp�&T�؄�����R����i�5Î��z[Ԉ�ɼȣc��^�Vĝ�\��-��@l^��ibܚ��N%n1�`6�1�������D��#��ka�[&]�'�Q�7#��:��)�6 �^�?Ō:��AJ3���@�K`��Q�����U�hl�CEd=�-� ���~B�m��lb/��=v���	�Fnu��:�^QO��vR�㩅�1�8�5�[��O0�f��o?����+��z�`4Q:���D��h�tqOW��F�l��E�d��.����J 8�$]�=OҚg��T�������j�ɋD��Uq:!�ކ��x��+du�`�����H��I�Y�d��?�����L����Q�B��NB���+�� �GhL�����YwR�[�l/](�μ�b��J�V&��{+��eÈ�&'���������Oo���]�)|�]ƻ��4���*|Zl&�ٖ٭R櫾�P;�T}�%rQyV,��Z%p�ݍ����əa_d��˫���ɐ��w���� �.�#_y>i������LF��z��l�7ɇ��ϬZl+]�����<���Asrj ^⫾'�l�C�.���zPX�Ԗ&#tV�d� +5�:�*l� �I7O���,�h�۱4W���,KX��� �.���|����t̥4�\�T��?�S+狒瘜a~?�{;��˕�ɖ�X_���K�ܒ�rуTH�903]��!�G�I&Y?��
�����X�k��]��`����;0�����:��N)9�<L��@�-�~�S�Dح�f��������h��b�ߊ�%��~y���*��P��E-��V�4��&�$�s7��:<���@�����C�G���F
�n�RE?x���;C_ۊʩ�<�ۮ�o.!���s�Ƚ&�1�&�}B�_�*�8m��Ϥ�����L?ǂ�e����fK-9��.#�\�0xQIbD<�x�w�x��3�� �X3Q%Cw`x@+k�qI�~��[�YD�k�B&m�ԧ�G�#�(�I$(���x�;�5�1$�S�U�P���CxP,��"�,i@��ov���W*p�����~�1��@OB���������޷�'��
��а9M]
�%nxn:"=+T
D�ңH�DJ������r�s�ƴ)�{�i*U��r#�:�"��V0j��ৠ���e�Fۻ%��i񼗖k
E;[Yh8��^�O��!a|�\�~�j6U�
$����)��o�K&��uk�d�8����_)��k'��v�:T����DVK�*q ����]�-G�Fb�I��1-� \��ú�"��nk�=����4z��	2���#�?�n�#��PU	5�lX� x��4��Z��E�1���.*O���;HÌ�]O�a6��b\�iā��n/l/���ެN�Q�j}$��\�`a�������P\��=���tE;�ؠ�/�A�n^���/K����#,���G���2�0��1�����:��Vis����;�]fo��� �
��G���� �_=��R�鲯X��!��6�w�Jo�Ğ0�2#��������P�g�;�^-������` '�.��bmUA�E���=re��nW�t�8���aC12��L#oUA߃0���4m\��(�/W�yO�j��=EF�MzP�5N�p� ����*�E#�Ǒ`�z.o`A��("�C�/N�����tѵ������&�+V�C5��b�/���^��/�ߢqjl�v�u�Wo�3a�u��"�}�"y]R50h�E��(�q��`\�w4Ν%_����%�t�>q�4M����	�RTV��2C�v�U�k�f�t�B%�$
SD��r�Gy�`���ՇY`*�U��ڸ�+�e��.���"�v��i�k�zQ~.1��T�T�,�n�G��N4��֒�/�{켺}�6���?�x���F6i%p�Nj���������y?��nL���Յ8�{q�~���{!��C���4	>��\]G��� ��_���G�A��n����}�<���A&�+��3.�'�IR� ����`�j#wZ\ ����L�i���g�m�w�{�Y���K�Y����enA)'=�lС��������,���>'�T�Z���-��ԙǿWn�0�Z�H�%|���>;��O^���V��Ց!��
�o\�<�䇡o���ȧ<�:%��m,N�J���@�w�8}VԖ���87ۦa�!�_�4�J0OSCX���4E�P�jt�Ԩk�M�u��#w]�fƗ9�}}U4Č����?������|9᳥�K����CF��Ϭ��=>ɭ>�AL��:��s��)Xp���^�S盡�F0NR��~�PS)�v?Ż��B��E-���T�j�]J�d	)��B���:�'�-�y����ꜳ������o�k?t(��3y��;P�v��+I+I�Ԁȧ�T��Z8�nE�^���E�8r_���R��d��j:? �%s��d�f�9�B?/|�S$㷶�?ٹ;%����ذ6��Ң��s�O�����A�� &�z���W�p$�X7i[���]U�qJ%�F�����8��p����7��B�弽_[	��y���`�uc5�E�_�7S@�a��D�SG�h}@C�1�h�ȓ[rRz}�)�9ޤt<hRf�S�ꛬ�~������ �q_�- 9�{
��A$�OZ�(��"�^~�*��i�w�K��8���zۢ�5�L����g����I�/�b�C�x�z��<�iz�"���3��(.���ɘ	���[J]v��.O�3�➦r�<��:���fV6���۶���)���Qj�$�1G��e�D�����U^߶�,��U�y ���8�)N5�����[��,�Ns��¼�U7 l�ٚڱ@"mI��,=�}u�����kd[��j�n�ZK��k`��f�pH=���#��,uJ|�.e����W?|�T�º�&u��:����O�[=�-�f�~
��j?��n�WyP
�.�HG�6]��DG!�rV�Q�9��}YD����[�q_�|�H�ݏ�O��ԡ�BS�H&�Ӳ�hB`���h�5dm�b��.��_�&���=�?��\�[���Wl��-�I���'j�f5�.ǶR@�"L����S2u�z�4ʅ1e�#Hk�%2�aT���&&��t�7��B����l�.V�Cn�{���.v��U�r�Kݥ:�C%e�+Z ��|,�ȟ��	�3��*��D����d���VT�Z$O͵���|�P�d#��\e��k�v���m�}�4��f��
��\i�?�l޾�y�9�DoL����?2���> �B�]���}o�u���[ n)����j`�l�ecq���@�p�:��ef#�d���\)|V�ݵ"t�����H��i	6�'�]_��'�љ��6+Șm��,���L�ۚ��ܽ@�����qei�)z����<�]FT�Hb)�2��$�g9ޱ�����B��l��3�<�#R-BK	-���C}ZRj���Ј�ؑǗ��K�ԣ�c��X���x;.�(k��FIK�{�&4���oE�5$�!G�M���2V��[�ڎ]Ӭ��MOJ�2�a���\iL�3kDf���;<�`��d�1�݉�?05����p�{A�n,O�UKr<��QS��*w#�JӠ{��I��M�;VL��O �\���UeNrt_�y�(F��'!������#7����Fn��W.�Gm|K��R6uGp/Z�R���J��Dk)+&��>*k��V���]_&0���Y���;L��ϕR[�ѷt��������Cf�1xɅ��ӝM�$��C��<�[�P��}�P���v�^B��|K��Q���<Q���N��ؒ^�+IGp+t	 �GE�o�"�9X�)`18�	8��3���y��g�k�>H�WE
�אn)�ES�xь��t��F�sX����"t��-�G"	l��`W��M믋�c�8�MQ��"}��6�-�?I��,&��0�xȢ��)�MFNnW�_�1��H�O<��ʻ���f��t�6��Ǟ��֫/p~��"ȇ�����lW�݃:�����-s��q�9u���`ʝ��s��"0}�f'��ث����zö�=n �J�{��Bܘ���S(Xފ�����A�SU�`cf��uЪ�Z�����#�2���3�g]&��u��}@��������e6l^�<�["l�/�=����9h�7�� �"cNЊ�)P��)O��0=1��$S�ߩ���}��j�g)�XSt֍��8���-u���Ҫ����i�m���v�:�uQO��G>�W��3"���%ϱ},#�8$§�Ca�w�:IR��7��/�l�1��xE�
��s0��p<r�D�dl3�ΦxǱ��?������Z8�T΂���$'WQV4f�Z��gJ��x�CLヴ�=�1�9c�9���y׃� ��z�%�d�{�3���g��_CSa"�u�q�X�z��R���
�<��ۗXU3�.��G6�>2xTW��!+ʕI=��ŗ��Zk�{ȂW�Ϗ-&����$�/DB�,Tk���qv�J�J���V�bϩ���hE^Bu>u��^nKsh�644���,>2�@L�Xk�L��4Sy�a��Y�-�G�����y�ށU��`�3-G?��|'�۴��~�=v���2��O9��
x����n�v�^�;�mj�#����I���E���(<�� �[�m�� �V�`�%|���AD�Μ3�O���#QM�b5-�J`)<�'R�����m�!���]���,M�X����PpD�8���H��B9X|#����P�/V�O��'�\~p�hHfM�?���V1�2�4RVj�9�yn��~ӄҭ
������1�Zc�,_�o��[�l]<�bC彎�&�>T���Y]��>O_���-�Ϳ��'�;x�N����7����F�5�uR.���j@f�\��
��޽[��f9�r�W��_Olk�;�����b�����E7�����ؗ�|[.�7Z�-lP\��E�:��l���N������ IJ��cWy��_�y\��ʊ�`|�f�Q�9!i�J�� �`�DY���